--
--Written by GowinSynthesis
--Product Version "GowinSynthesis V1.9.8 Education"
--Fri Jun 10 14:53:22 2022

--Source file index table:
--file0 "\D:/Gowin/Gowin_V1.9.8_Education/IDE/ipcore/gowin_empu_gw1ns4/data/gowin_empu.v"
--file1 "\D:/Gowin/Gowin_V1.9.8_Education/IDE/ipcore/gowin_empu_gw1ns4/data/gowin_empu_top.v"
`protect begin_protected
`protect version="2.0"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2021-01",key_method="rsa"
`protect key_block
YNu8g+Xq82dxlN9DEXhHt+1Uhi/IaQOaAdIHI49LcWG9GUx0xWhfHIruQ1m+gH2qr1FNjk64Ckhz
GNHAsTG8sUyb29Sb7OJx1jNoyiw+1OHhDWXs3d2KqM86CuGEXZmjS0UaRe9dn3v0T7lTdjCOV4LY
sTNeW70AC09fw9k4phnuMm4nMND29IRhYvrtmhx2qCLyipBAdjY0J+0nagp2wvrpELTL2bxX+032
MjAxYV7rMsgJ2yeQiL31QsBAgrVPEm+pb84/xSU4Inj6hXmuyjha11zEUicLvKKq+LtimoeMeJEV
+w1DIunDcY9+PEZ02JrMRZNzpIXML9O2vAn25g==

`protect encoding=(enctype="base64", line_length=76, bytes=97072)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
Fdorie7zNLTeDHCxEi4NCcELqaUZP5NDhiEBH2vtNbo8Oj9G9ez4wkGF4pJi0fPVR+DfciWEu/bM
Et87rng8W8lrxStI9j6pscw+BbT3C43LFsZEl2WVCL79NeG98zyZ+4sCVsu2ZjWXrACO8Bt7DO6D
3AgpiwXfm2/Mph4xxPyUbqCGjccNp4Bc+Bi8wUQ9/gbmxSI2f9JML0EdklKa0jYHQBYfOaO5DZfL
onXuew/k3/B28qzFjEoQcT9u/fTVgAqZYn8CyCRh5TiNYBVakQnnSFJZEDkUirmKVszIUywYMjBN
cpepdUDP+TMLpICaQL8Fh9nnbOWDTng6r3U2c/C9ygnMNldJ3jO+J4aP2toA+l7KjPKILWXPVyEW
Z5AIAUEByXaJ3np0TYZwZhVHpfHtCUa1b+03krYmD9uMrgLoOCRg1PVOghzAM2bn5AEPokQBjq1/
HUQs3kBRkGmPmop65fvFOPbWRP16brcLC5ToylPe34THy4bClTsAMcTDVOuQRYNGkz8yjvs/qhgt
XeA7PVmMFg+ro2YVq9Gp6Ebx+B3faWPS+88HACT7RwbAXuZsPBoeGphzRJwTbFVTBLSb6wyHA75z
t0RVe7j379wUsqLCPXjqaQqVt/8Hxp5PT0+7fRy927mR+VhZbwUPCqfSRfJxyO28MWLZSxbQfbug
rDEOwsi5yrXAfrtyqBmJ8r8qkvQzsTwCczBa3gwY8cQoNDKaxLBDXrfnC0bY4hu+YD0QMrSClMLf
nONq7kyL2+9Y7+XrW4jk0qfZNTrcmY4aaWsZrLRWvuc81QKSdwhy3EMu2MduMF1AyJ/8LewKja8L
DgDBFP4Jd7cC+6XuqfAlpQS/zK6vAghE494wZw41UYtNuAQieyLf4sYpYIlFr5+0yasuyUZj8Tw/
lxpQ/ArsKCwZWU8KH03uNnziPHS8R2TWq7ar8aD0Gm2ncjAYjFkJRQSFM6Pe/85GhnWkdAY7q8Ni
tm/hPsIi1IcK+DXzsLvM8s319SVgsGFswH2tsVvXn+OoL4fK0myIy8Zhf5PSIPcsOctZavDEB/H/
vzmzGD+d5lvCe3oiIg0paracL0qqiTl9bQPzUertEUpOV5Qg9zJ0pRoIw0jyyQSGoSR9+CpsmDgL
xDT9ZS5xP3yGAa7y5KHfW1ERvIo1CYsvccRbAgpREvdogCDJR2hj9jweVzotGpeRLcAWzUeu8npO
z2NxTcf0roZAalxuptr0aAUxx5z1nSV2MiliRTX+YmATt/zK/8pQvpwFyBr3oeHm/eAGdRok+bvs
cnXMVGD7ovAVg6YS3+XSxFAWiwdbjYS/W7WOU/481hO/EidC+gVZyLP88CEXQZOj0IsoqPg7vr46
BjkUUifjhVi89UCg7IXvb2yNScAeCBGxoss/V4Lx0VEy5Ab6E7sICSvrYjEAbV5p9F/amMtjryq8
q1Wyp+X59RvjkYEfAP2d0bMWKEdnBQYO84bsfXtv+Hz0K0fccy2BtnzD/oN414JTRSapUu75jqu+
BLYJN2QwCrxRjmGLvIohLDIfEer0GbxmEa3Ip9mfZJsouzgCwBI/w2aa5TOSGDE8vDFQ1sihpuht
exJO2ntcO1RwkrMtSeyczsgPiHZlseDP/2iFTtttdu3Q4ht9maHgpxWg7GiEN4lqeNg1jAHZhAVN
DAw1MZ4bKXd5ylcP8Jp9NNnGUddNnOeLWq37GpQlL0wfIwpJZDDgQM9F+jF0dvdk3tLgvhU5lb4e
pBjOIAlnNSRK2UDt904hi9TGuuIb92ujQ5rrzquQG1MY/0ZOpniHIuKYkv768shr5cQOlhMV8QrT
Z0QaQTJsg6D5JKlay5hoQhJrUGlkGbIKItkqhfq1x/WGu6BYbSyv/9/yErKwWnC4lZwXfQ44/Wym
piiR02kM+wwGy6mpvattA+1vUWGe5s3q89EsLfsXUx/QRy2cEQorxwPSPs3+RKFyO4srRF8Y86jH
UVsmfNIO8NuDQa8ItKNesauNtHayQZPLajTSlhPzWSYLw8MDwnYaTJ5f8Cewc1wQn85qcpUnQvGY
ZEOv5F8acW5//48LNW+MQnGtueNgxt+g8dSgWfIbr7KJYcagk8UGY57quXPmk/+nNkZC9a44M8yB
Bc1s/Rj550Gcs2nZpWIlSLhnvNumE6UKfD/uDbKsqUO+tuKRnivzR4pP0gGvt05rvymtw1h4rVQx
WuQTcyMew4HkJZGAuz0JPL1KPnniXDMSbHmk5QAr4miyaY13trVeaHFTNeFwUBgxSW9AoCd9Di8D
8JBYpcO07CIVdW32wgAnitWCn60s7K5ls/8MxpdjN+7GUW2EYTcZmh2AgmIIA1zuQz+Lk0lL1avz
5Nu9pToo0uHc7Oa5bFDd8cd2xR1ztDD/OvTdssmbVtfGteA9J5Y4sxr1u5UY5f4Kb7D4bY8AEy7r
IpY2hNBVSM+t8sVIhm3md+KAYvUTG7TbLH9o3ZCMdAhmMxH5slgay0nDEOgsdAD+QzZOWIdK+EbM
QCcYS8Emap+IBCJjqGtQLejkIGEV3xrnHt0qRHmBM1wO30ntKwMo2uIkuWiRWg6vDZBGEoF68hPn
waWQX0NXsUbA78maWlAqlAq5v7OLBAmnwjnY/2/nGd/HS6kErYZQ/9sC5+cVKh70Bb88QF4QGH+y
2e32+N0niJf900wNnOcrxhVwpA+pdGjGFqiuk7WLnGsL1Oxmo7FvFyCNLQakz08mizhKAmehDV2e
ZT97p8RgRRqv2xWjjYYRlgF/Op+Vz1PiATAVSsVGMB7stLM4IdilK1tS2YQR/Vp9Gffl82Vf33lH
jdXnoZYS4QY3KNSimvqZrX7DPh2cFzY3BX6epqWPzdPyhkTyTcQ60/49PfCk+flkjv+7TkRifRUQ
VAZGpYxJXjXagtzn/LtcuHuCuek9Apz2sJ/amQt1/KA+vr9Pt7b+lWNnUZYSORpFMny+tyik9WD4
JrI7cbpC79t6wA5HPTDkCn/88WSds6XQobBqCK4Ql3Ti45A/gki+7BnCNOq5MbnCy6JOszEgyHh3
/F9UZDq/E0BXe8gdBcO0j4wW1BqXFGiIbvaJSjbG2j870kiJ00Vz1Sb0F5Yv0nZeaViXw9bxZGFe
j0k0/J0R1HNmEtsz21kdLzB44hzVMeTWO79XR3jh79iPiGjh7sy4+076P0oMLdt/+/j0dpGmKL9q
lO3HttoonwncxxUsvwmqVESNtnwsmU/YbOKeMTW5WwM+qwwHBvfCH1m502vaAdLZvk7+1wTNioxI
2kKCaKNKN+a7QJ6pHjsBmFGq6pcKGAHSHfdARK5kod2dFogz/BIALHgeaGH0CyPwbhw2O51f+HaC
2a7y6fN0xaAOF1bpADUlf7eWhxkxJd8pPFZgFZw3FsFf4fOE4dwue2mFL57/lny+h7E1K6y4cJUH
Weccs4Re8xMQJvXnW3lMnx7X23u0gjfyTrFeh4Sc9r4qcx52e5kRqbmFL1dhl1WXwo/h15yAYjgJ
/0R38jadZZBGwKSN8vRwIaUT7ZdZOaCdTmYv7e2arQjxgtxrKxN40CSArltbTQKRVv4hEsypgsnH
2Ex118a8FZGP7EIUhj/quCc/IFuscSPdNadH1IWUKX9wmutgqxDvGjwjf4TeWhaWn2LGnyjAz9Xu
fyK+pdytkK/jRtkIwt3dC+i7GiZx8FtnsdZCOzqadObYx81aVn3eAnT8dkL/9wPRadOn/cJDAqg/
pcCgf9+8x8+CL9KSMI0TBylA9iwhWs0QtnEOV51qIgiUBuOBzcGRI5PXbXubNrugkhRB3Vz1JzMV
kBD8goGjPjFPf4y8UwGjg8oWIPr/n34mKE2icb7y6r7KMuoE3PxzXWklsg8IyFDcraYzFd4HVzhp
pmtQmVaU5bYl3bLxNpcuDwkNHQBsGgiM0GqjECRWdRp8DKySHxbExfA/Vra61ZOKtH+E8drXrBnq
LiZAqcN9T/iFEB2NH+0EgsmxhSrK9jq9idr4jzuur91/xQXkzSj1CcKWDzSvx3Mp7zBngkq4RtV7
KLAkHdq2se9F5jwxW9lYhVjtEa7yY1GPzE5YiuaRJcjVhcoqTlrQfz+VDFwlcW0p/WKDwFBbvwWy
TolkSC4VVHMZNe5nzd+ODWa18/KFETviNsgKmShg09s+8K6znBwAhVS55Yr+26NEHnrDqo6SNLBS
kgbjbLRtjFYfTp1HTJXYvpImQbETthWv5v5dRo/I7NwtqGKLGhHBcOpcRM/OR30NYOdyvL8aTMYj
6Y8JpsNnEaAorxrcRbNxuw+IUf3ejadz97Hi/p5ZQZM/YpEgnOZgfnHuGa85s0Im4B+lizdyjJkV
N31/Zf/61J2JlWph8cYlbLGnifMjgJepcgAtTNcMfnINpAIPU1lg6cNRVmgxY9BfsV6+RvHNAdHB
Q6/6KaQZwEpbe6lcvLG+QEZWEWBl8udugSUspJeRIOscG3JjI/oqxxfRLU+2fzLNWWJap5Ruz+0m
oHkAEhxBuDDTkdODKYh6ieslBu3W/skDGkGTgXirXH5ia1b0Z+WM/56+bVTNH86NAp/k9gG0+J5i
vtJ6fDxDIkuCzGj5nf9kGXRA7d7SlS1a00qcJ03QeolxZ4yZCHlkg9buyBIOBJ3aVR7wYbY1Q7wd
qnI27eAPnYRLoHF3IzQYz8RWVyK+F6IT5H/h+WA0BwcdGGeEch1DNzN7UjhijINpwCKOTJQzwr3Q
ZPjvkWm+1HmaxawGiPPJM+pDv0Y5lF6NrvYcCECvj+xywlT0glOHNIRsO2CC7GG3w51k5bMmJ4Pb
iAyifohRNLtsw7jzzodXe/4foTWwazL21jnRhwjFwlP3tFyztfa2Vn4usuqnmdJ1zEl3xx8oMmJa
7khUlmHDjofnasVPIt1i8EQjPk83by6cJ1IHipqDzfDgNS0tyxQaq2pxIrBJ+Kv9AfQpnx9eqRiL
yLcqZA71+fyL/Jtt61667nn1em+uwK4yRRkeXj3Sr5VS2pIVONfEmcUKSUK+C+nWlhJoYCmi7Z6Y
rmH8lngmDMImBVu8ioA21e1gBnuOozsMo71lGofu5e1jMOmyOurALu21acoxqfLH3NlzRUg/o33J
uKe1O+eSduWbq8ukjGaRKXez4i8u3sIFITi6jq3vOsnPTGVZEMdrXjq4Ksrjuzs4aIZmLncGudaI
X5ePW2/k5Tze3QRH+UrhJltezwfNX+Yi77OkMT2DN3sARXb2v9hq1q/hXivGdGiPskGLherjxguh
Ifk31yY402DzL/179Xzm5xNg5UazRGrxypnXhUO2bjvXv7PsCipgQ+3OlQ1aCMVRulWhHECFjHbm
KREOeKs+BcOJUF/CZyzEhEuRvV8p/q3r4cwpnZiHXRUBwuJqc/uTT3UPFobuCJNbNF5h6TXXYIK7
NG/WAl8QaUFZeFTDVj9B0lgJDRg2KJ8TqdNMX4CsV7zk0idbCJaoPKtPVYlUT+J8ZxetNR4edVKw
AKuYxXgjVL+JSFh7G7HLwRPj7M/vZylxROdPjlBuFhWes3Pg7k5SW30C6UyagJEgGb0CbNVWm1l+
BpxhfsIXfRj/7VHsW5jYeLbZ48YjcmnHG4qDO789tMXMkor43LtxF1AfwKaEiZWpKDELKMsT5pJk
VgP/FmPUCRUuLUnUcC4tN4g/krSUyjtIRC3mPAvKCwHh7OAdaZs7d+ZYKw8mbpTOt0NS8PxJMRiK
ek3CtkI+gRXFh2++28bXN7Q9dmzXSXlmIKRiB4rGc2/gmno+Rft89YaXrvx61uKhSe0Dk2dm/EMx
xjzjY+gxm8GjlcUKRrdzscWERoOOLfk7SJON/Y11LcPrkKvEB3MowK5mOJPKP2PEFKttvyFGsTVT
dP68x93x41CQIwX3oSSem9hEJqCNdd1VNKI5dprmVkCcwdFoTKABV8dM3LU4U2eTqwUv/VKCOBIl
El0Y4zbrIL4sukasezrM/xuumR5N8XodiNVrgqsxWaC1wPX7mPWM+cB99v7I/fkW9V5lzl8h5Bjx
bKxjaCcdwFitQoR7pcqlCdb8/uF8nXUOC5mgTfiKRA+8FRlSH7nJMcTEK+7AAyCcre/Bv+G8NUPc
iT8YDn0cqxjlqZEJu2I9m2CEPxlb//H6FAdn1qU4h81d2e4WaLyFrCRGumKuTriPQF59//3YzRyT
qgWe5GV1KakfEcVQuBHF2M7Rh6Rj7/MHZoWc81JbjX9RSQHlybM2G4qS8npEXC7OheyPcB/TiKEU
5PSxcXPqqpOqp7IIhYznrurb8s+2SOWtCw06gPCDWsRxxIyfIFy5epntRr2SlviaIl3lX2ijQK7A
vpwqtEO39X5qAdL0KDGIQ9x1/aH9tGPebJSk+3sUdnd5fiQVWtd/8QTgBE5HZZrO1sjU2Tb8L3Vd
QqORKJnJr3r9COx+xPtx2nVzvey2EOVi1dehr95yLGzOg4+0WobY70t+BfyvA84XEVI4TS25uUh4
9dZiKJDQARietDPKbSmFnD9FKIttKYhzWJWcHEgXD3UmIofoOOdHeinwUbwadLQbbSx1eOz/DwQe
RosqmqvtkK2PQdM9OtMVg5l3MVygzhwLmYArhxD8B6LpRr2uqRkBdfef0cjnVq76KWyMVTqc6ZNn
ptkwHPAV+yg2FeT37+ZA8R0v/5Ylzfn+A8T/PsXYQXTKnq2pOMXcSWXJxK+OiCcr9AHKSCWo3MOb
qKxKcRLoy2ELLrs6iJ+qKXnJNFZG04lX6bOVIpBPJnBF7SDYYCWV6LHQlHZuLzlyY6ahZouVOOmp
k+n61qMl6kxyWPDMdU5dHv3BfShXntQFQDiLoNU7w/aPqxt+cTtGrrDTJWBhSk/s2RjRaCI0YVMl
+rprn4IWbydNyYxjOpEzPHLCAyE66kC0/M8wa3/zTGByWs81fehitvKLRjeF7+KREVhBjwg49M9F
kmlLnjvpGCp490RRAdyotQb8WTnG/M2g2Q1MySEEvYcqE6NOo4p86okbQC9TsZxbM2+xT5yVmDTl
6BvESqEDz3CRkgyQFf1SXUzJhIxtALxL7rzgaIlgsdlBoCWX3lzwIeCo4wXm4ZVNA4ytgTzqCGVW
MNdAjvhxyMKGDgR9od7Ka/xalyXuB02/L3yUl4vaG4pNDOzgyWIKaqHC18IDs9IgwRewXtPZYcoG
ClTNNxPbxS+hRZJz9DR9Qyo/OaI6wCXRNztyTpL1pkYnnjwvJrcFRkHw7FBMxWjpnyZ1amV71NgP
24zlva5hngft5YKtCqh/PY6ySU/PYtjnkpJwCI/A2My+0Ro97B8II6ui3dzLbJASf6mlwtrmGA/1
NgfoNL4544FGX2cf8012YJJcQ2dLsV6wq1vxphHzew398Ir+jN8AfAG+qm4gCUNbZ8a3fxOd5Tft
F8BeXgDlcx5j2Jn+LGUPeWfKxhKsQu5lGamPuum3hw7RoQ9z9tQ9Z44ZyTrepSwwxRO7hxqDZJMU
eYA1o6/vYt1wAtkfMfpND+a4gspnENE1T7pgSxXKhsA1NV9hfDdqNtYDuVtTLG1Nvv0t9JwJzokV
bwHz+9ctbs1l8O8J8aAKSQTM6chQy/7nn3UOMSowLRl5Z0xtw2FEhtz/Dc/2/Id0qeczdZFVJfHJ
GEJJ0YxFMakNG85pbKouHagVb1Sy2Iz6qIp89ADotXZDMACxZaEjAELUA6mmvNgLe1fD2UheJ0aK
5GJp6lQYFaGopp3P4Yz2r/tSj6uXsTZ5wIJJRm0pWnq4fCEtIReKnDJ7XEdSdSaN+iL1w3iz94Fs
gVFGmWLUgPIdaK9loTjI5qRY2yeWsoT4jA8tB4qw9yUTcnmZU+DosNlFo/jiNxptlNNfw3DmKxaD
afuaG4ePKfMHcYo8E8eX1OtJ8YxrLNYgvNcPt1GIjtMRZ7uuYx0tstW5Vd1nPNsm7ExtS0kd9mEp
EdoyqWws2OTq+Nl6GZRpmmMNI2Jxj+LliBDInKpHHVpHctkboMPujjDpOF4a87M/2EySDH1nLoM7
jB2Qh81ppfGPBl4GX2ZbFkIdiIiYRNPtq4P0zVtrCb05kBlx5qh8CNOiXIG4jAc24U4IipGECaNL
NKPrn+erizfQyGFnI/q04gIQTFHyv8tavt79ArTLhVlxMmAETO1fX02WxgPHgOZgVtj0Fr3yFopy
5L6RHxXn1kpHt/YXLV6HAasV6iOzKuW6fydrKKK7NJ1IB37e0ORwj1qNyIgcxHbuCi67Z8nPJeXk
ASFfNSXavfckghVY9jiNZ/lmaaxIEbuLp6mpZwpGhzEjeTavhjQV0lsiszXnbUkBtA9XB07XG0+W
3Me+jGbQMlC/NKn3RbBkpLes1xvbRujoJoMSrU3ayV4SnPe0+5v4NwA92RGqGJzDdSla0wFW28IH
Dvrtcruzlr/6+XvVzGjKH6HWCCzuBqri9ZbladEUTbFlSFBlnZB9uHaUguuqFm6sfG+i7VY40g+Q
c6Zw0P3Ljw+oebuW4zGrUSPQMWcGfLQzjjDakBnVhJrhZnGNZRGY3iupzNOLQxmh5gCQoPfXTwuh
3h8cRqsHIy4GzxcmSk7P0hXW4sS3bgcDCdBFBxa+uE8gJNacV0/bdkRAFv3PYMOdBkZ+cmNBba14
DlJ3utZNLBtkv5Peop4f5og7Fy57lN1GNDWpjZI3U1xNS16yNdI72eRcjxopWOco+VTQmimgl6Hl
eYey1u3etGxU4KRqLVvQeJsvcxfL2+fdpWxXV37SWBTUMVDVDSp3xFK/zznibGz0+4lzxHME9Tch
z6S4yyinqgLwXMCAH+b5VRxmzTVzytPG0ZJoSXDtRfgJpUyqpoaa984wqZpr8sKd+2DQ4DhBHLWS
mYnfdfGCwZOiR0Y8tde27uyElY/6ZOLXYDUpmQu7/WpwmFNPv8KMX0BQIXxq6FBUN4e6C1s04USx
hU/BzlfCIr/0XeR3ZMWEBq2Cl3UmoDBsafG/GqkPB7EemkY6QpsTVDdpDroKbRo/PmbpduyYflBY
zpASEPzQk4mO+xmcFSg8MYwt/Gjc59QiQVJ/pFRG6Z/zyvt8GEfD4CEp3U3HX8MFkQamAL9grbf+
xwwG6tv2VLjbVfL21M7Lu7n1xE1Xe3niB/RMOMK5D8xqA52CC9N2wI+J3qWpVL0x1sPxN/gDJJqb
twk7hWdOTYJUmSIHgil2EO/nYkBj07m1od6yhOrcAhDrDz9PJc9BbU6OoQ8PmQa/cp+uXuyvrmuW
wUojl8dA3LS+nt0QlFv2fTNVm9PlE/w9mMBN9piqg4z1Kdt+lyEfccQjLs1XI3Q+j29YhLafoIa1
HcV5304RXn4sQSjAwcbzpNDwF2SvqzpLxS0pGI+4ONWCVKZME7hDzdV6EPk5Oskddf+r2OurARZN
/QcmWsI3p39SFuMJVDD0SH1Dafs8UZkIbgdRMF+5B6j6rUc6KcfeHCipuwVwi8GTfNFjOoHPdKEW
omENj0nvBsVYL1it18G10Tl8lGPILg2canPLO7WZW6dlzJf/VTYzEwGaxCZEj8hTkY8UGy8yURNP
iyuk3Z8h5El/GiHyQmuV46PBlnDMwrTL8Hysxdjcbyum1JeJs0WHGlFedMbbllxPCn9JIvRU3eSS
F1uBkcZs8ESKJaE7I/qLjow7xVW0/vw2thajfdD/1LoMs9OXnxfY8WErDmwDvAjl6KpsbzRcjcAt
L8OwlFbu64WMdpqSIBFm9WHktBHu9xAbKx3D7JC7aZ8QY2NgO4I7RYdH54yH65pnLJY5nDdoziKe
lY9ICvOgPen3F8FfBe8beiPKbSFBEcpaNnDBI7nsCYucScU2WlnaCyVtx+fAqY4fwtHXlX6U5tGe
0dHH6LcqHWgCBcbno5AscFTIEJ+IsAPsCwypPVaIaM9tJB4jfLFPpXfPH8wAUKJB5twClPg6wb2y
V7CbkICV52SSGOi9okBBmlmZfvDl2F3Z+OR6uDxaEZ2otYhCzayKE0ie1GUlt6wGFeoMMPjTbEIr
QRuQbMuhAAqV4vzBsHRd71vln9Tj+pRskl7iqb9nScRL6BxJyr4GmpMCRus6Bb3ix4MwhFteGHuF
bD3FHWqvNmWOHsxPBUD894QdZmys7dSL3IY5a0K6gTGJGzBJ5QgLtYv2DCuU1rapvdNivcbjT8fE
3RZnoWhp03IlO+OSFOFquDkh8hkMyjywmz+IfK5kVwQZ9CXWDOWELA4tukyidZK3L+GgssnCbAVs
Mh20eId0P7js4/c7nYFAvvjxHYSOgnDBvujbzIGrJsrmW58ZemQ9HDSZWXtr5WRyRnLJ9X8XjA9K
TqLpDrwuE4mKYKkwFjdjn3F12FhVks1xc/ujoO6S4ZOq0Vbzp6tlaYeCjuGlJUr5X1TqTJu1f46H
yNspJD16Ec+dqTzoJG4NhJzzPWDVTEIXKI+6ZqZGmdsOwpu10Q/9ET1sOIN1iDDjMH5nrhHRDjZE
EBjkElm+Si66ZLH/DBJ6QVaTgoNBwqKNkmx1tZJvaCCaoLcJCrVzxtGrmd1asuK6CM1jZynaNG6H
fslULbt4S6cw8KRDUreW3fXTu3Tuxovr5ix4Dj3lOLkO4GmN2PFpjRwRH8r+7y9l9Upn/ExW2FwL
rOu0lFlB3nZ8Ya9rmVXAy2ghBZyRl/aNlwf7PgcN4GFUM6i7wmQrO30iINVaILqKizdSP3g8Jy4J
gLc7Rs3CEMeHMG3v15j4fSh6Fsbk/CQj1eh48Fujoo4dJDnTMma0SAfzEzh63oXB8uN5JMyapgJ9
iwhwsqoIOyEwmkZhAJiv0UjUuxg6ESL5iHfrvH6yxkm8Y8ujpe+6ts0M2POXAGnamnB29sv0WfyP
O8mJCS585MTp0Zf9qKnW/kZx8jcVxt3t6KGtNcN01Fy5rAB+174gL6euYKxg8My3/QwhrCXjTIgo
E/3aFUhyMkfWszIYM6I7IFNUbMUjp80o0Kb22Ei2FR32XjcEndd+Q3s8PfK3dlF1m7JZC7qWG/zd
fzrL9heajMiz/hCXOtQ79xXv7stVrijPZjfKQSlPMtxqU2aQtnsMkqbpUt50cR1xA3VYsWV6LrtG
3o8vmw3KAIxDOYcoh3ICpiT+Ow8wqenTP2tv81vwh6y1d5cR7E4xP6vsDUHAVri7JoQFGAGb/Aqs
aC0WAmlwDnLjvHWl6QFhbpyPwjDi9O32xpASGmrYiACdpjVusx8aLt1UCggdi70N6i0ca9IzFhIn
2oV5+ymRX0tindu++27/oDfFXAJvzsyBvkPq+Jwl+/gBNPs5MDA6I6vTlPC1FuBMHi8sYfmJxtKx
DCNCiCeEtxgbq2dKDt9MtYyAdpHnMRT5VxgJkQ+jNwVZ2fRcNX5oT/R4LOx3Y5NiG/HAy6h5H8EV
xNsmAjmbH/p5+FyopSlhcsE4SLlAdMa8tPaWUfq2392QY5WNzlE9s03eyoYzizzmLWneOrymu47O
V5T3X1A3K+Upud22K/JnjWM1ZqMKADxvc1eqzIicXMjXiMKnYXQe8rFq1JzhN+KhmDOZjebvEM8D
GY8P+Ao3ZRRojse95ANM5GwVaUyvrkOnVx7zEu0lvaC6NaAITkxJQMhRWcLWbWdQkI+lDX44L/KD
217hXZfvPtlUecjFutuQeUjMDtdWT6JAohjNAljkcnx8qG7ctAyTekD9i+9gMkOzxpW9RUVeinR3
hqlZLFrTmt1khcOh9ymOJnOxvIhoBBgMKD+8hYjtq5wemYbbDRCn0I0bicrsIGtCgON8tK1mbpST
jdjOvHTmlfKYujl6tw38TnlrBPL6WxNj8tpcTmmQDFO8CEfaEdMw6exvOgNXqyXY4ZFvyHSWZkQM
ThJ0bm+tscz9PmFDwx+kSGkCEcA5hEYLI72rYJmXvIJPfZ6+MgyNPe9oCvozetfb1Vo1TOs70/n7
S1Ox/gYkY9WVTWQGIJNX6leeIiHnLGmMpJ/1Y3U0M8AN5cXLeNoqK697tFBsD8PGMyS0ZvIsbq7M
I+KL++h0wfKu9KV0Dezn//PSQxMNqezgcjfLbhL+ZAeZGVvHaCMQZvCKVjZXjljJj3WGdTII/XIC
YmThhQtg4EabbJXejQnIp9855g7NNwk9/Sp62OWGGLjz5RpaIRgfnztVupeu5tV5KVU2COBJge6x
MAGWJLs+7JML1QhPfumylP/NAjOACrNdI12ztq59VIFk3LSyVfGgxIBR+fskwHOxsuXo4R91yO8B
90dweTQG9068atal4Wt9GWTNHGnZ+qtXFv7HEoYDskLyJUk4bqYv1vwOokkw8RBMFZMcT0jih3th
F2T84Mn8rv7sofhu4AInIHmrUj7+MLL7zx+g2YZNWGOrPwzz4y2LNBsKi7gKqiqon0AiHqDVu9HO
2RzGPZ4CMzVEkoSRdfjENyDWPmXp4c7F3eR+srtpRUrFID9pJOWU0mJYjLGBXOMuOVlqKLzi4AdF
n3rBHbBVOCcWGFQU75ItlXQPshn2v0M6SN+yk2h954k1krEUF+xHjcKe3MmpWuEhX3FNKbI5AOhq
hIGzzG+aaXj5QcaHwsDnBag7WRnvdPNgCnqAxu3tKFhJBVV+sqm6cnHOxDcU/sH126IHg6U2Ia05
qJ3JXFVeZA3YbjlPeGTAYfrLGhOTGBLEaxTTYlWoO2H+UBrpIPrSp7f+HPy5s6D3rKJ/PAeM+ahi
A+71jZGeq1CDZpPsHIGy2fzMnDLeaSxVw65ax8hDmhtyomEiyFYSDe+r4v0caXNc1A+C8VcRGh9C
Wf3NT5TSsXbPzPLlmttmCCr499sxRTLfg+CB8nbcTABvNi0YTLYeHNGqbJZ0J7ywRQ1Q3pFLPuFv
l64Wc9o4MfzTv6NSI5jHzV62EVc/xy6jZP9gZiZd/nUhkwkuJa065s0/AbdCg0ZvTCf4KyT0ky95
r1t2yW5d80sasmmXMceY21EQGuvMJf9mP63uMMIVWmHqK3xLUXfSOdGztVucMh9SPh2QnFGLPyzh
JcMvzD1AEl8Q3g3YvJwbXFs8xI34yt6Ksv3xuoUGO4Fh2P4+WTVd6h53gsiweXxn09Bso02UneYP
cym/5w5QjwaMOAWPKRZqGCrBqUtt6JA1cFtyMc9GqKjHbPkaq6OK1pydtER3Xl+Sp3+kbQk749YF
gTBucbacQeisrNQf5CX8VdlI8rrY7b56F6HZBOVJnnERb5V1bTn5/LOhb897f0wDwcujvebi1Muw
ojCQcIhAKr0J2VU1MJfM3E2Nz1TmPIjAE53P+BDTRWlJVVfxcJMx8mF2GQkV+h+QnD+XTHwtehdS
8W4Fy9bL9z23gchQAnujZKe2nuSOLlI60dpTlM0D5eHWa7JMu2pkZNGM30Kdw5M8MDZ0DJ1O+nGh
L4PeNlvV+axQHHLBaIyVWbkEr4g6syO4485ENmVol9ox5o2BEQS65qylEYKrwink9NYA/tsLNI16
EJZDOuSf00DvM95Mnz1zojMG7eqq1etUxHmScV38TDM8Dvr0AeHZMApKt45uKA6A1ikJf5v5NMat
eA4ZzAKptKFtJY+ogHzvO/s9qLkm/T6nDGRKMQ5vi72c7wN5JPWp5covQiuZBGUrFdEG3Nc8MYdv
X/W0tzGebfkMdA4Ytm/FNZBbrKaMpMJPfXuZuEAqC32UcssLXD+5r2DTcqrghrmuXrLQZ/pmgb6f
C3h1aunpH3KVjESem4KroGAVyQDE3IOlye0vGM9sJvLj2N9Nnkk1JQnRT6VC8iw6BMND+UElSCZ7
9Ri1JGWJOw/tMvCQ0zzSCCUwJD6CaHi0mDHNhvX8ZQva//KYSfwgxrqZe2nyy+Ffi0yQecyPDJ7l
8Xbil5CAc7AjmVkf+h2E7fsaoeqJNjGWWrkBGiVjVDNnPTc6jsD/LaEddVm8CEcSxsqBTHSt9zxc
R6B2+fy96Zm77r2d8Ql+wCX8A1taDNEyuJG+84SXQ9UcYKFD3eaKlbq9EtrVJyzEumV5uXARJnuw
9pQ1u1AdItAZC51sVe9eVwf/H13djX4Upb3JnS+Jflp6cE6c1a+ZDfctaTrVkXXLLbs7ZzX25FXM
RK5ZEyzD7gwZpNcU5nUqUfmlgKUw0Zb/nD2mVCcLWl8d+va0omrfVP8T8wKGzqlVFMr8njfdJ2A5
cW30d6KP+ivqwm6G4zwg7ASUN1sZ2AwLnZcpLVpck9NS4Q9soJTdTeiJK1Q9BAWJDBQPIdrj5BvE
E9CDCUVuiWDPuDpt9tnsAsDZU7dmlGPzMvVLGpxU85atkBTpVYqBaI0DXCZ20utMRyxSbdDjIBps
VM8rEVxIxR/63I+boMYYDYROHhdtGG8MmWD++Hz502yKIvsNua8DWaSE5g213qE+G+/NictFnVbZ
w8+K6cbhlWlui331yktU6JcxP4IBvNlUFoBMlH1OC+7/nZesIWkMhF/wOEy27T9XJ96veZjeSvEw
1jBKux0cwzqRUzIV3724/cjNSnTcTBFUJsbYkKf6Suq89tTn46Pd2aLp8QNzu7n0booWPTwv2zQ0
GD6MISSmgHvijQlgFPR6Rghb86plWW8C6Np8xGsajiKta9ezYogETjKR2k7bYclDcq/AEE97yqUn
emou5571V1645WITzQ/ViAh2mQMu4JC0zaeDk7aJCSkrjp/H6cr0LUIPnvOh+UcZ9BTTpzkXpImb
6kqO0gB2gCqC9Pcp90I9gZjkyXok8mn0uAG6HHJ70zz0csVTLIFGdm/c9npvOOp4svtP2u/4KKJr
j07QsRH2xh+8BfT0ox6OQ9lEYnv/X6Am7+fhs2PT3dytxrq4S8IjTRUlbpW0QPuAOo0FwW+QxCfH
44E23Oo2kku9xbcrwJKU+Y3k3lGa0aPgxTNqtAfkgmNrL5ZeJFnhNB5tfCusCj9EDok8laPvBMgb
rei9tDaJbDD33Ga2KfGePCiyOHS30XLDvyks3/ZJqzL2F1IT3VfxF8mnMbuCTGxJLNfacfwtyhz+
tcaYDaTYNbxHbbH6qA00y5Ktossx1SK5Nt4T+ggmzkNLfVHsmVgyY59tix2e7e5yQ7janNOsYMCe
IdH983WCoQ9977gYBEj3w6PAuJkQq1KgI63zUbxbjvurlajf6BNEL4/bkpK9q2JEG7AVZU5fI+XX
zpCUqPNhV7y1a3S87QOPPOCMeSNdpvDDSSf8ZFdYO/UnHAkZyNK6DkdkaPstXVRg4lB+iWYk3Qtd
yy++Zihytj41HrFoVU4PDWb7aYwJxfziahwWGdu+84HKOXceODjuBtJ0I4jNDmKnC3/Xk8nySZLD
R3NJRY/XrUWEqATie3OsTym4jID/RiTfZlNTqeGLXrOFzVRJ5MOZXXXKLmomlNV93YaUhIr2oHRi
ywpcx9WcKNdGqopTjZ11og1JBlqhgswHc4MIxOFT5s48D3ZQf0S7iWTeKEgnQusRr2JJNLXHi1ci
+0qGty/DMg9dHlgWGQFLl+6Cph6CuMVoHYQ/5laYFGtTY422X0C5fTc0kpiZLfVqHgUpBCtZZYe7
4X1Ug9VmDFak9zEBZqT94tDK1Mmj61qjCeO0cm2JqFv+lMKayRsYXndImV5cx0gbn5Z0hhUUBJka
+F36Or0ubbhEv76l6+XcAbFo/SuvY+zPHyG7VxOn/35X7bPGM4TYYaUCgS8OMCbw2y4dfSTitlKV
rhKDFIICeMZbv2EZgv8hhFI9gjvLd1PQqg9Lvz0i098xKmXCEWuvfFTcYojLKd91ajMJbugirMnW
hBQWgSXXFfGnPkDxIygdGEHxxEocLogY0wa4XPWt592GRq83Vfd3WuVqY8EO4sKAemCI3Nql7tdF
sFK0I8gJc302gp8Jvy60oZhOghi0KgesNYVAYvdQWglFg7DBvGX5bMTCdCcKeJHADuTtupGUxxVm
Fn+A9OWzWW8zA222u+Qdn8RBcYfzaX2j7JKknsV6XJ30fQqPJA84y8aH63Q+P3HZkrB7ssMgezR/
0FumvnYrVdI7Z6R1p45fHdQzpyI6/4EQyAdiDy4FnoKIfr+4b59HmN5yrd4eVaZdzB7wiArczUzQ
zVqNCLSeXnG2HOfX/BV0lfFBlFtPnOH7SjI8vkNfJ/648s9hFYICGs7eqqQDU+g9k9mEPwi+L7el
l41jn2yJ4qxabWYI1OuizZ8nCCoCav2pv54Ij/Q6CSQJ1AnGw+HYepf0u443/QYSLbIFRug7YWLA
hfLliE8ljWr9OKQEFs44oZk0u8qavkXGf44yGXQb62KOrJdzP+OQG4rDuolm1wEZkvtx8vAX4mTf
2DhGqA0II9hkn6yr3GQL7emy4w349G4uKxMvimAfC7kXeplDD0bT5AlAXXkht7OEsBepTKnxhEJt
4xnnuQy2F7RzBW5yIiujY0FH+Zc8R/sBqVmUK3iDc9GS9nwwgproYXSnxzR8eriDuszZgemwmbUV
PllP+a4nFdudYxo8k9IZb16os9GoI3KiT0Ag1V6WRbCXZQ4soBqRlftZxV0YFXFrtoYC8JgFCBek
ueB+yiTv7Uhy8dlvhAXaI5iM6eW3y7QwmZucy+JpTR1zfUemmQv3XGbdDPkOaiyjCxqyMKorz/LY
gviEz171pbMVQ8wY+v8sEAa1qonCOPIlI8HZgkizuvy/KzIdV69gmWxkGem+zMudOyg5v47xRxcK
AvHS/Rlv+IZZ7ljsX8Svu9bU56LIbUzyYucCMdm19Epb1KIIOtMftvZnTc+bebhh0+YGcoE1yFlN
bFDY3mr5al6IOLYapSouRXYvXm/vXtgoaE07veCdWaPkrrpQVcyqmBvBlmPmZ9AQyAnOsNSSsNnd
sxOdGmNpp42+a5ANfe6wCjfdhboIoJ6cUxQDD4H9nGr0PkOK6/FDKuFi6iGKC+pbualoOWp5wRZO
RYV6ZxPIG5jtfGqRq0/3Bt6jgcvoDc1UDA9nzEIvCf74dXhAbS+gaLbeScVYnUVth1cHgAGmA/Zd
w2rpxnOFnphBE4c3zJOofK5wxGvK0uATNpBj9SNSN4OuA9KuQBq04H3Ym9zO1g/ri0u6p/HifVF9
RkchTMqvzH5jL7s6HdjG6V01PobiJ6C998juY1jA7IQw5vnQUCy2+MhJ3J130q1KtO8y0UNTUOrD
SDgIz4Rw1ss/I/nZ0g3kjHjPXImpGHHnre5CperIxm51Yis/lvRqknUABXf8FflEWbxy7skHwZxW
Clm0a/LfMBIHTp5kwIqpTEJ+Ylx4eyBrDQlUYK17yEwRTRFrGQgHkCjVdZq7KClLUgk262k9xjpu
QLMgHtMicQ3LW9MsWmjwMYJj0uJb9zGyd1jtRfu6UB4f6fvPZobye1nw8W7nWUdE5Hr5IAzNY1h4
sls0wrY8prQg0t6OoTLdNKShHq7BshYt5XwZnJyS3hZ0JEsRukSpsrgrUC4NsfOBRQ+rVExfFjRz
bLksbgNrjuoJ0BGCj+i/9e/WF0U9tn9VNHrmT3WspRIPdUNwLGtF0HsLIKLAbV0DTyprOe361hAE
phQX6EQiHL86i0OVLweVF5UpyyRpnbSLfz75aXLlGhCCg11r8RkANSqgY6+TW0i9UupRlNmJ1W0J
9UZ/e3ybvgwKDz8CHd+c1YiMRXz72e8Yam9/QtfLBmiAyWeP1JHTfWoAar0bKcZG71MrjnGnwsLF
SfoidyR86YXWhbi4CVf1LhUK2N25hgp8TsEx9p1iX4hLV3Qsdiq3/axi19zUCN2CWkxG7h3eqnyS
gDoF0B4gx+9iO5iTs7nAMUmi/wcrr6XQEF/sJkrIKsMyG2PTZ0I5aqSDToDoC/TneNIxXHNZIE/+
4Tdrgj7ExNLYf1UM0FBHk1IZLpPRFbEWV6GY6xhWX6fBAVJVY7HWbFpxSnOItGIjLMM9FcPytuAt
oInedc2sTAz2ko1/4xE66Nn9PoWP8taodESuH8U8RDduKm6pfVEqbrz6qNn7ZL2oUFyLnQvbKdf8
wi0AwgKmcaNjNQhnYhkS1leBrgNyTJ7W/OIaKLgZ8kfVHNpffGFKDh016O9cHCocKK15fmFVnxkR
ct5ELj/5XgpxkTQvipvVZC8bSEOxPXdz9wB8U3uHHbiJuUOdfw1HZsSFOSVHMK5WoF/93gXn9VRk
buRYZfv7U4DMqANg1RTGbp6k7yMqLRFVCAeuOKk3bXkhFULkkihrPjiHcvvI2eHF1XN/spPhU04V
4FxplAGyW6kfne4hmgFVjY9WiQaUjzBrCCOYKIhU05Ej6qqDsiAxXGLEgNRxFMZON1Mp0NU3CsOh
FrKbWNDhx4n8VTzBCke+K8dIRaxnVgpNrXNU+tjb3HlR1+ZWnnu7NzdzHMLl5hBU14tcTsOgVqwU
1+yFvVJcLvL+V/K6RwTkBrW7meyGyIn6RX2NAOUaHwjXwDuZXNDWmRoBcL5/eDHzC6FjCpiZ0ggI
jwI8YylrlFoEQ9PMgU3JHXFYuHFj2xGV8MBEFxuWbZB9XKcmDTTzSIfPeP1N91Or2kpD71llhmNq
p/tOt3U9lAlaxlECrRPfDP2iXcwgYMk58oT62U7XP4gMeCVCK7wtDNi42o/7fN02uPxJkUBuLx0Z
xdNEfnfnUVoKcVidQJ4pgDXZyuPYwNLlFkwr6ohiLMkrH+gvrPfhJN4k155K189oVr/zOWqW2Gfq
pL+J4uSOPxXlk+YtdayNc2ydHadPME3bau06or2nz5ZjOcTQ5rYXDV+1mBSCEB+wfC16kVIFa8ag
Y4ndx0Bp+SORnO+yyLQOFViHOo/kAW0ZrshgoSE8zGodpkvD5zvVkOWSPHUS09iwge/IU4iDTHRD
yxF5Y51yfHOqn1cr0mnLl1Ai/LawcmCr5xICEboUk/FOT3pv06FKmJ6JNFkwKSd3MWR9nrhyUDWg
YkFlWLTmnXkp6AyMYHMkZA4tBvTkmLIMtBYeOCPYRJglwJACzDysyivXpdtSK7fLQDP36wLUyQf3
hsZwxGp1nqIavAqq6qG21cwlt2r75eKfjM5NzTCwNzn1HikhsH1OWiqZd8r2EY3Oi0I/enKNAFcG
Fj9FP3NMq3Tvur1RFtesY986svwi0oUIJjaTVCIAy0SHz9356tWDvsaAexvYhctk92ozCESDg8n0
/rp/6EcdM/QNOjOjoeMnL4VFsI5P72YJWE3OTN822f611X+R4qGKkVWqM2PD9IqO+9zziqO32ooz
LGSUErqg8pqNhAWhTFMPKA3GkXznhszu38EuSqSHRzfRWxe+dvjFWNo47zmBi5bNF5KiZcyfTGh3
nMZ3YRzsbJQx1+kQ2rCn2PZAMAjM2CBTSXroB1Lzi5gQgv568x9jdZoMHzZu3ICc6kY2gG2ZWj55
RcqF/QonEWS2f//+EkBIuE8PGXEalEvKyGEgNjIaRIwsI0dIxeNANXvj3Qr20fdB2hRkhE38Thib
VYuMJbJ25HgG5E/JTUNmDEZ20pZtZy71Pe5YC5NF+y/OUYjFUt56qSFR74KOzlxWqGwfjQT8SNfu
sgE3a6zK4apE/+hq9b/gpm7jgv1XITidIDvT0rTqucawarCgcGWMmxhz71kbqt65RTKZgn9Ive0h
Uov3rRA0/cgIALcE7wIkyKn+LMMt8ZzauKEEIZz7R7zQY6jFdLr+FiA3cLcPtJ5tKWc/OkzCdQbT
mWWma6EyXWplceZFTkNDNunRqdil1RzB2Sif6Dz9V++UqmsWRSpjKKUe0m0qj+kP9z5ETuDEhBE4
UIywczF+utDCBPjSCmUA2ZcStnMuSsddRacOsJhxdDTSGSEOYsFTaMc4PNUBMh0e2LDyeGDUO0XK
e9u5xujtXglPKWS8qnSgSO3lp63Mb26kdt/Wu0HVYa5v02xKMBzNmMG0T6SewooHKZxSO1W8HeGI
B5TNSEtxxEOZovdVHYYIWD5F22up5Iza/xsrqSlihc0K2QYr6nz8P5xMRU5ptqYxC5N8znHeTISR
AtVfume9vQ1Qt9v81z8OJlQhfT8JHSfCVc2SCB765n4oqq15CHgAS1lBEVKbQDLvF6rU2z1O5rLm
cUOK7RcoYcRzm9o+WHrwUzAy9bMQHQnNwEv+32d9uMFu+HTWvMr/E/iGbg5MXqiHHI4T5BS7gXMJ
93haX7JDtcX0BrCsuQGr/XUJ2hJu2aKlQYa41wCs+QMAIUAbPwbWYJZL5fqSMhf2GR759rzAjd00
S/8GnHS7Yi39GaKXq35fJFP5LrADh+ssI5ZddMesrPYJ1MUgWBC6QXcV7Mp8zLoZ1kJjltCHJXRv
Aiuu5Xy0AuoHJ4sPq2gVsH6E4Eur1NsLFBUjwX32W6I7UjGHV0mJrPsFpKSYgdV/7vH/6UZd7j/b
o1XLnRl6B6+bwCrzvWdzm3aAduBSqCbHBjSC/VVtv2VL3aMSDuf7QbmMxkIw51hgWUfbX6+pxOVX
kyHFQ6u5e67P3tnheF111pgg5c+E3tV0onS9hrIxajCUojYUPNfrUm5q7kXaf6FeRiJwnLx25jFi
pDfNrNsMmBx96JoprdUb8ti+ua9TFCg8uuok739Y/vZW52Pj+0gNnG3vkdpiBrDhmBVOHmVmQhnm
NjuiFASPrwnW+PZUZoX4dD0bS1f3jBk5Qu4wtkm0WPpdSUBwi7zNyiv/lrWS++Xh1hX1Fg7cTTvx
q4FZSRqrSNQ/R2vI1OYw9n4QGX9ZpybJQTfdCGDHvpF8v2HH9tr9QvCAjidzny6qgn6+XJv+yciX
OV+OffNA7lX/DvbrS0uAn5/M6Fb002v6NBjq22K5/yGol2Z1tnh6jf2bMsrfQ1TBoHBaDOgOzz5R
9JHfNgI4q9y1MR82OM2hCW4dHTO/FmOAlnLQMcl7IR6QQWvhLSSE5ZPcBXktSEJnCaHJP5j5yBt6
gMWFKdD2WzmtD6620wHxdjQ5bE/ZZbI3DfE3t6TcJsP7xldTqgXcEsC5h32tPUcl6t/Ca0ho70XY
eat1zunaeXC0szly/4eAvuzp6CXAQwg7F5Q7SgUKKwXgv05C2CXbomJ/M1VWoH1yJIOQLb2QRexr
0zyEdcdUtTjhw1QG/SpzdXnKEoXOciCBMo5PlMfkkSbH7inNlym+pcG+ygDKUhY6A3xObVTGuNaq
cv7aZcU9ixfko3wio4OVXGQxk6bONMblBLLykKybvHZ9eNaL5eMIUrdLD8Ae+izCCHpTM9Bx7YPd
PrnYEsdVVY1KOao5QyVAPKIf6Jd/adVPZbYU/Q/hDKMJKPpMVfqDnGpE8oQzqQbrUrB/EUY5yICK
is81skni2cYq2gIFrRefKnSumC1S2uFr/F9u6kR70ybzviEClPbEP8Moinb6SsG/cA0vW9lWpte6
m4oa2sPeHLyBYD8qWU9HvUUJbfLEl2DhBlAtazKxH20HS4Dr3RH3HEYxp3wHawCIsZAWsQIqeK7C
S+kvx/PbvW/pqPABEG49awGAVwakdL3/L9gcTmBh1NZv8zxp9kUB826G73S4b2IaolxIxS08ZEOm
lo/C34Cs2EyDKdhknK6rexGVKaFkgr09YclmgTjnUgknOKhwGaO/7wtk4pmAbfDInpqAWPgiC01p
dnEpEQmSYZVCr2/ZPB1IX7rbVstFAg/aZcXFEGA1fyDKMALDExod6NRejulxFwTrV55omP5huylU
1/JBhflMmz2c2TY7NqM9kAdG/nmiNFFAiZdokT6c69bHpEGxrlqqjzvc0YFBn5iqaa565xfaBL5p
D376r8GOyuocurWLYWwlo6PUqcdoQsv7oC3SkamIpuvuWEd8yyMb47BksNhPWnO+VMZVoCM6GWgz
l8ZVyt5srPX2/yaYIstg577WdDmYpXvrZoPf3DgbZaVBykuQQhKp22G7ckRpqTI3iRnmu4GX9T2a
61O1YaCjvhb7/mhdypiFjX9IxgJauJhVuUXy6IqnOl6isxDGAjJy2OintEeCrOSp+H4WVDmz//eJ
N1+rYU7G2mB4yErMv0qHHNwMfCJvmI+E/fJvv2ydI4mEtQuuKnDYwxt8ukxUIi0lj/SyZ2j9WzYx
E30beTsA7/lg+7/h/ShAC8uJKx3i9NHcpTtu/z2XHN2shC13LMdziXrGNZ4EvLF4KiK9eP5SX1Ge
fKkRZDAdoNaZyKdm2kzm1EnrVpbhMz24TEu9GK83qP6cjSw69fjv0oHa1z+k4oE/TBHTrK2ZATVE
qGJsCPdA5M2CQDh268RjgDWAtRuPCZHp9wQJDAfCypSgWAasAxTJdtEmus1xLYBQF+XzCuF+VisL
omqbPnPZAQEn/G5JQ4FlKlkXW0TWy7ohgDm1bFBNbcw9sDC1TB7N3fSLvC2lfwg+G74vumMh1LBm
VkGs8Rh1IrlgbsRAd63V27of8glEp3u1G6R2lCFmgMTxYY4h43o+4m6tLs3sA4rBByz4tt1S952T
s/D9SPsBq/zV4X/ymSX0Uac8RdPXxEjF9tOhr2z0bFmtwaJ2WCq9eyKqgN6AqUzh9g0YqdmzJbTv
vLuDh8EyKSs5cPdxtq2cktXYUsyi+JzPsRvGy2WPpvckjrkKdNNCVmx9e++zj5No+xsDVvgza3Zb
hOkP3ak41JjnMoSGhZPU5J0AH3UIHZUXaAIFfmBx4I1GZCcClPDtw83ABv7JB19Ftbm7wkn+wmxd
iICLH2InxnS11lYCK3djJNc8toigcnmMQ1Kdjx7FuQ7eFXRA4t4fRTrOyPPvBArHsmOyhUwBuf3x
SyrDmHzRuh76g2bmyAOMrs7UMohOpR/Lhv5nRLxIuNdtzvPoLC5xfM7cdNJHQG7/akb2vLGRWos3
via2hLkND0XOHKk2zcKv8fjZ76I/WVSGiebNM27V07D5szgnhFukJxjHs69wA55UO/IUTRYdbMLM
g6GGYZK3AyVbdqVJrI42PSavmXcst/YuhnzubL0WGp1RShD2/rQanJTXOH+xyRryuAadnXrQV9RI
NDWpR9+F/GVEHJ2hTq00FhFPSvCw8seA6iOzUAyZmwtN6BFeoh0/mv7BeLSgXdAr76GKLgwi+QMu
fg9WOs4ea/7niWh5QsHaG8MHcVtyL1kgdojOxswhUq7LJ3RxSoxlKp1IoPmb1c04kFVMjWWqGDt+
WxDimccy6bimbdRmIOWoOuSDvX3P+5VPVdr9cPbLuCLLQzh5pX74wAxyewHw/I2tTuabflTsNc/x
zAzw/RdlBRxPFjae6NL3p8fjJSo10LGPo/Fd7hthr0ukJIDAHwcxOk/6c9Xf52VmiSJuU0urVsUN
LudBGQjB+JisTGAvjWY+vj+CKCnl+HN4qu5FE/vSi1njpu7WLmo5iqCcGY1jO2g/WeXXt95Y43cq
khcfZgU4HjwATNfMuS2FGfg4BPRuDTNvR0hF5UmwiB0+lvzhvelSRB/9tN0gY+v21a5QewfrMFZQ
q12f80piJMJsZqtAkZbsbWcPXTox0CJb5rWFXM837VypInceUkPZSz8ba7J2H5c5xixn81vW21o4
v7RvL6tuRXqzFYlxELiKPWu6pmG+Am3AobxKSrGPugHBfvL7gkuoYuejfR5NNNjHVWZgf0ZF4daS
6n0aQ8bgCOJe936mSjPG32oBeowZQgIKLo7Mz1W9G438WEhx8SHvpjQzZJQDQzeS4vQ30OsxD3sj
pF6wdnfDgXVN/aUV4k+jhyNuxhnAoEKt2o90JKklcAushtIwxNTUuVacBdgI630pFUrzVcyCYZ3Y
4ZKJsWK1KMyWGTJt7e1nvh3JSjuJ7P7DBcYhOZCROojk4QDYUli1Hj46Xdw7m9wq7ZTogw+bbBeK
m0s7/eYxGXFtykYm4WC9GzAQf1MSwkBERdNmu+Xa2d4atNB5FkEZDbHv9OUbE8Oka5HraNt7+s/g
7DEdM7zRbyhS79VALNcJ++l4cGTL5WMiTe84sVXYStvGAjAz6XDXzxynuGRhVgQ47qk1xxcyvFyg
b9YR3iXBLGJttByh2uNH5sRJmmpOZPWtzYT9M9zzHDST3QgOUmZd9X9ktb2jbCcXMjeC3kZUIkjp
C7o2ZKZIInMNctIhTx5am3kX15/GI3xSNhe/QVTZklaIdiESGoddVpqvtuZqFPPAclcWbNrFU5tC
IZClZFIv5zB/5UqQW5XklxaKQsugTRjjMO0Tv71GHiD/vT5oBZC5rRkEQxfXOUSGeMK9jX1n3ARL
aaK4E+zMVR1eMRAlWsm4il/0V8jrznL57PK3B9YOak6N5kdZ4ted8epr0mKUChiV6FX2t8aZzf/j
63OgEaKMzLMtjplgehqkzUyduJAJx+0MaSNZUtt5yetWwWWL9aGKDy8zsmG9uetRXiB+/0rK4WqT
MFGr2T9Au3sGi261214TENdxIYM1e6iyJ4u77W1Hojwi8Q257YXMo13OugNHVTUURcD1C5bQwLU1
8J1iEp75eOQaHzyam8RJAC0dsUdURS0Y1Kgjy0PzT2Cqirq8C1Rz+eSoqrZW5sdmNvxLajwwzBaF
BTisiSd15GGtKaydaexzHMHqcAbq+3OArXT0olu24r9fnRIQMRmEZS1TBom+kcb/LD7XlL2BLNFt
kqudpZgj4s4AXgW9M77lXghnQqb+qChiyzgLjeadqFCrm43I/yPhieUDurD/nyJaw8j1zkV/d7vW
BKkTlMrh3TtVwKhEWNAzhejGkmL1N6WN0gtHu3yilqsL8xajxWupZpOJtorNcr9PVSGYG9Wm+1kT
AVWUY5QiN4PxrmJL+WKH+Cuvr1WRkYEPwzEw+lnpGufYXz6Bts8lCyKlQt4NQ/HMn/eHXQwE7UDF
a+UiRCz/lUR3CoinNH8GpCyX7I6DT6gdStdn2rsCdt9moK8LhAuARcRMwmSIPXbyFNaUX3CXM8/4
miBS+1CmUWCIuD2kuYv5qE353w3C47D5GYvryyXjnJ40zx7byrXn20iW8UCb+UEiLO1CYjMB2y54
nKcKDDmVJZrss+TBNhBXWOwV042ZayRb3+QmHQJctEJvVqCxx+xLezf+k3dmm6LEuFweK38EBUlI
3ZIXAMa70XIjvBT6vJBQWpQ2ZIB2AtaYInCoatwttbUcbBGingM/+tG2oQKAeAJ/OESF3KGm6eKZ
LROFDreU3hRZHmwvUwWabqH385eMB1NyjCcaGKBEEFsxr2XXO3egxQv0YxUma/1P47bZG5vIGSNT
oJ0z45AV6RQt56QrEyKRITxvtKZyZTEgU8aUgTQPYzmiqq/XvIs0Dx1V07y33t1VQh5NTq6L7eMJ
hyXsPDK15XHiuNHtvc9dCChq2cIQm19/Cb2e8rXkEByFwpb7j2PPNXw+LUsmtziXJL5p1f0kGk0+
3gQ+bqGaj5N06N+ZPnW0TClcpzvCIAAq0kFdQ9ameFA20YU4q5EwW9LwHtpLe2wElE6RDM68/JyG
kbIiBQiAVU4sABH8yC2DKw8awzg8tnk7T73VbBk1S5qM7zW++rNve50D+5IT+Wu9ly/cBxAUFM9J
NckQ3A31xtrN64W1KcKidqZH5Ij8DF9vJJgMw6G5CBMoTw/QyubvjdQbb0zuTAR2Sfc0qCGr5a+S
/tHAvo5q9Ndn/8tUhEaQpZ8oqzlSrvNuVXssxutQQGAH/h54LtdTLmTtMUPAiYrh7lb0U5hu8Uck
iwULbrnrKEvetTLHMtafA7D+ybm7t6/WDQRjV78h8nroomRoYJFO/qX7MRMA1IdNyWhAc7Crs/cR
LuvdQYncv24CJsAYgxxl+ARn2q4CSdha75Hu3/obBppeaDKd8kL9vVflYlUteBYmkyq85oiy9swc
pRcDt0pCjLQ5karSaoGKI2NE0jtmtf5aCDayqhhgmRt6kyO8P037lwVLvkzmcdFLb/lSexEzGiWM
GB84cPOPsSAFyJ/aSGuCYdTkTUSsQdiJl7TQDxHlLfWolDhyFsu+j3fZSyMcfKNW+iQoSjaHGBUW
vkwITIzbmbHROSRXFtukZkvfnJ7YAhzQHsmaTtaTIbudSaW1T5OWVfAAAV584Jtu+ps4WB/nzmgD
qJdp+EisRXy5r8FPecKKKsWZYO90kfoyD1NFx3Qm9YFXQ/m//EPO7EnsGQXMHJP3c3yx56ud96Mv
SPJz5j7SXZn5n59Z78KdWEk3htJQTyKfRUr5OC4c7O4+ojDgQ4YJfXRkd1JU06EvJI8ymmjff0e7
8QloVC1/jpDq0xm6ahIF23lMVWmSfZvdQXmOSSJ6/kBETofKAp6DDf69PBRBwg4gK/81j4jABQuv
Y9J0vH+o2YRiZdApy3uy/khhJ1hgIpKhPfQCg4dfe9u4LTZub5u0yudYbaLpXVKpKp16cXqBxIsR
o1VRvhzjn75Rn8S0Hd3mx4Py31NXshBh/fs01uOjIRmeoDcOrOTNsK9ZqPlOimaJi+xuvdamSshG
CFbKJaurI6qAadJ7OnQ7Nr+TSm2lZhabmadXMwbqtmTu83mjV3fXtBlmGSmOD11uHbtVVhbZG2vP
ycLpiyfIW/dBlvTaBUthTEClXvsgohtakiXR8qgSBpvK6p/F1riFap3Gk/asgR9TB0iiWkuFizAX
g0z2fzQkv7zxJkXZy91m5nwBIr0EHhwowmlVTYe3pCDznVpViINMAXRIOyLMrQhBP0y2ncx5N3wl
HFdlvkCrjpz3Z9tlZpdPJOqJfvVW8NvdnJrQkgJ3okwvWrzLn/0vMvEqY+uCTUSMiNUO4qb3v2mN
0831jTmhab8gzVldLC1TpXa4yQb1orb9q7h8K+U6SDBQd9jb133eHrYu1fRjiLqahK5cHFzTaOGj
nUXADkC0R4LRVRzLeW6uaG0ASF8LGVM9WC66/0K9YxTnwYaNwORyfvEHqLW45zsWIHxzPphIVd7N
rRxugCvfbSgGmdcvQn1OE7RVrkEsnKKDYCTuuKp4DleJaHlSvE8bRdGlEZXuEjTf8O6Io+L8lrt+
IzNHKQvfZYx7qHieHNgQrQRx8QDfw0fkew2LDfJ8xXLnWEpHWGm1TfEhsEc2YGtC9sJikrA3MCNu
bznNm6Ky8yv86IAKcW8mdtuTfOuDQgjcmoen+k/WTxOQhovEyYX4wN2QkRc3/WdQBNEYDqw2cox5
11HvpFX7KaiCiRYN+APTOjgkvKh2+TRgMIPNo3xUGPDInIa819rFLSTXG9TZMQ168etZ3eIxriNL
9dj5dbZx5f+JA5sGkR7p1a4uvj+yCxn5n7+2LfuRleFnsQqoYwcYHE3p15VcCOkY7LoPriTUIEQE
J7nJJyF98rqPAGqdV1Fk/WuMXsQLI7wAompUkxIv6F8CMRiaqtuPoJ0SZJ7rJJsV/SuPbPHjWa5U
5bBQYZ2r8NPQf2QWljywdJfb7/kOniYpY4IdfuovmtBll/OXRdTcqFBhpLbAt5MkAzqq488K+OOi
Ce1TfUuB5nfLqZQpLTEKmuQ6YX3fXLACaZq8LN7JkppJkb4ckTpqnEvtugNpTlrnzTvPmXdodSqr
kP+e5xM3ApI81EMrp9m8PXKLfwmhchUnoMZiDex4PmLZNxTr16Zk44eDyP0nVgA61ZUxxh7cvvdw
f+eY2XxYK+2Ad8STiJdi/A+s+0ycCtmTxlm+x4BfrIhFG8ASS1ojwRcN8VBi+1g5GqN75eq+XjP0
eE5b08ue9UdzPp6otAeJcWqaeqb5HYjNL82heVL2Wj6w7FiQX7X4kOAADARUgkY35z2/XRttMF33
pPuSBzc134yYYqeoIfiSuAYkY8+eF9zDFSSyfw4BBCGHTaL2OrzageB/0mhg3m+ZSfMeaVvsJBjC
GzgFhi+vmeGMN/DM4xn+MTiAbgotSGhyVbU2B4jYcMtmmPmwbQ6DUFugKLosjJYYU6crYoF4EXl3
A2yEj8IUifuQqt+P0Jcw2vPpSQru8WBWukyWOmTn8zY7mbRija6dNDseaWuYKkRAydEahMwoW8rL
8U/1EjxIMPw8oWHnqqexIeMlJ/oCyTayXnEXN4pNHPsBpf3ZCPhJMK4WRpLAIVIc+5MToZmzKeQH
Mwj6Mhe/2lD06Oa+EXYnjV18EJx74zq+wpCvUBeEkvAqrP9QVS4mZgmkjngF6ipebx9U6QEdcIlW
0fPbdQwRl1V83pwHUvUmIx5BG1+j7Rv/XOLpuxJYlSlK+lGAKK8S9594w1IxLg3rEqazZ2ZFyKK6
ztKdDdps0XU/AzI8GHnCNeIcspQ86cIxs1T4K0urcat0X8OPy1QnLk6RpDv1Whqh/077bPGa6Rd/
9tAs/HTPmZzVgPMhT84tlVyKbPWIvXkkh8T8sakvc8Ozc7ZTUoqKAZyDFmZ+tPaDo0dw6njvm0Oi
Jo7XzfrVemw3wVPcOn+wc10cyEoJ0BWlXYbdImjzajPORovNAfe9BEYgTgN0gUwk9+5+cUv5Asxq
C+fHZfuulbQ8GWcdHjRduFMo0rLNZ/FL9aGHCVNicqkvM5SlAC2EhdVcoFgn5VmcRyeGIMOLVuYR
zZGm8KCKx2V4lBqtIQJru8z5NVuDXIicETFM4JRNkITPN+TC4/TP8qVg7XJf4vQI3byqHTiujZDn
u/VKcOmzimTE9gyXKNd4qhSLW26RjhMDxtf4ucWNFTxO6RgMaErQJlTk+VN7w1F5zmB0/+idJFeK
hsuxWeFmU0vlIm/dGCofWrmSmbUdi9oNK5qsYSTsbkmhcJLboAjFBgct7WnR8xoHP3fBLo1soLQ4
l3CCaKmjR6nZvLvZzvX+nZbzUc/ihrp0ZZB3TAWs/w0y3WVBzudRDopGtDUa2OaGSLDYK3BzBmTN
N6RCYKHIP5EwojqoP1gHxLFNvA5I27Yc2bhK9+syMc3OeR9fohyJTcxFJVo+xxjJDhSlOKJi27gm
CQqLII1y4ySYbMXWsVeZN3+VRIoK2JJalP3okqC5gBreoDVeIXknlKmlC+Ze/95kfaxbHu2kwtOe
XNA0qMFww8ORj7fJBREfSo5O1aDlUH144yRGqf2Z5CXIlsJKZTC0beKgN4A0c7UXFuxlwAjd/ekO
5s0KRJigPy6XCaNs2vXcr2e/AwEwYb3+rRzgwdKIPDbBn0Gnb27mrg6d825Il/FzOo11vH5DS2Re
thjY0e5b/QrBGeLEpyIzB8gYSPLgTjZkvoywqudybGSRp4jzDKH9DDWpMk8Pu8HogFUjPdfCgcO+
UyU4bnvDwC0z8j12BuvMBFgazeLAGIa6m3FdafRh3sldq4RxBkYQ80mCYfEZ9E88WPiaJfLoiqdQ
T6Z4XDAwjU2HwzZBROzl3tdbee8p/bNtWIguXXXPMRcssGaTr02Pu5vz2uG1VYoeoAoIRCJERUhd
rU/iGTljXHB0dzyTOUZVwOM8wofZEtji1bJD4nYzroz8XIQDhnoRB9CpmOPOQ9IlbAYGC1yTGWbf
8jolcLBFmTUN6aNNBWKoZUnbqpyt9vholfvT4O9rnj5h3gEsRAM2+12bCCELfOVUEyX75o7EcL2N
IJ4OzNk34749Gxj6aAzbPMG27mf0mWRrr5TBNleta99E/2ObxbouUXqJJrbQVYz+acIp+pJGJ6ET
u8iUJ9T4QSXuj5UUzdMJSDAo7djDjGJ1Q9Q4BYsnHtMQS4ZL3JyX64TKmN8zy0xdZfXBX1Nw0Awt
ldNvTxx0hMJqQDP2pexp6Fd8rTTrmcNpxUFURQZ1GDqukZigJwrZmrS384LVP1lzvTMnWCEI3QSt
RcKCQC7uPr/akY/ZE/JkEqEAAJpiqSrdibnm1MprGLfpnT0hoXfG6f0hmX00B0Do69+qC3Cacuo4
OJIkWAtaHGNJLSL9yu0UeNB1Xq6JwUCR6UZfBQoZkxbleay3FzMiSdV3oRL4M4WnBvCB542z0sQm
/8nCA/BOh1xr2yww05H+oC2xrfgQc2znBQfb53FML/u+0/mpdLQ+1qMp0POgNgu0gNP20jvCucia
aulEa/toreRrfztRxJkH2aURlr+YvD+3QPQyqjqU+F7vZNNGlGwqggMGclp1/uBnBfJ/VDktHrRc
/ewhamub0U5JlEp3V8DWmhJutYuTfqdzXhzdZPDbHIxOuH4TyyGnegaftBDomb5t3rp2BMPWYCCN
tiqIrqK2wLFPevmI60j8a/9vpGF8GoWasPgSZH/14gt2crBvt9+ciCzuDdkOkfDS/cAgAFrOjyjv
wRVKoXdB9iQdE4x7mdzamwjXfiCbiRoBwerN6HhYKmqV7ezDmjQ29Dn30G1/jJpbUzSJCffbQkg9
JDdq/epCmbUb1v92cDBjenil+FezllxvfxQ9Hoz495fI0hFNnDC+SB+eVvg/31vQRXcgHLtQUX/Z
bWfT39U2f7t3WObMZLgWIPv5RNU8FI4hYdJanuFB5LYFM1gKG/E1GGkpI9LlvHEk+qwukmPpM6V2
BfAjczpZVHI7oRdWhMLlrqAZ8V+BOHrObOUojlK9g8nlgS4wW0wfBFAeaYNOgnbDV0XtyU4gXaeX
7WdZRlW6OgaOvfGBgu27Fz7JPI5gsUSNOMoBggJnG0blGjmmN7sWmphp53kEStDYJgUeW2mryJK2
D2FdX3ZT355QonTYCh7RhZPe8wPfOIY43FN5QTyo2xr3TRG6QvR4eGm89E8wntYl6tqGvRpEDxEN
TxIa9JhbkZKASjBoP1/YxCR+brSIDW1CWDSbegSj1nOKYxJ2AtpoBaSwxXCsQuZd+US5iutMzKXW
CuAYeZH09Q2oFJTRMsNbEnBqxCKpYGy0uskx+9jZr53NOM4asAZnZ33A16N78WaGkYvyKi/JPJDo
oUejJdR6v1XL0/PaCKu2w/YFCGIBuJCHbaECDqsM+z3UAGoiISZcw3MxKXXJ0wEh5wcXX4tD+kl5
5Zoc0dnIbFepgDA5V65hQdrCqvaSiT3fnCL6qJWfWEyrIvsqWS+YRRIy+xgKwRVnQV4gZd7SdZoJ
IfbytAw7kDmw4OOboxjSVUKWHXBbrUL43/p2JiqyA9Q1ExCPUPQnheN6kzMz8kwVGTTeOR4gnEbV
bL1G2La+vLarPGiY4PMBmT2O4vCGPS6KCQIm+aX06ybNe+plCdC6dkRzcPPlfICDhLxkdtSP4SgB
iXWaWC+7URIHYOf9VMxV6uIJbDG4KFrMOIM3zVCIsOtiS3gvNrJ6riZnH387m/htw77YfNyGZIUD
ktp2URQEmSGLcLBVqbFu/WRfNxFoV+UvkBtTYnfdim+z16mUxwsT6mi1teoe1EDg2N5qcTLZngow
Ga1TriLJmWhEHIBNBVPp4XXRt6aQBNskgOAdYGdFNCzccBOYlw2MsW3n5QCFfpbE5TGqr+EvYFTz
W2WUEiBRaog7rjIa5z8wDzDwwAE4QgrQS3xVKlOA3qLf4bB3ZgxZZA8SSBTfWWv2eQAgkn1sEC+s
VBGLMaoc3Wbea0RQzN6c32ZlLG8JakI/cmbjpPB4wGAfwvukNaelinpwmUrZqiqftTX6BLXwP12X
o/7TiiGfKX4XtNm9BrQVnst3RrKHNEahUWuE1pVAknC2RZnfSqN//FRbHEgCU//aWRHhC7Jsw0++
tgq9oYP1mlLoKjsgy0Ae85B+MXaE0pwx6QCqSCz3GOa9XKb5cTYsUiXFeQA0Z2u2JCphnARCkRu8
o8YYhK5sTOPmkeDtibRDckS4TLqHSuDFn7gWLCvNe7Yyrd8rble7l0irZret2QTl70WGUMMG/eDV
mffgg/Rya2UEIxJIc/48Rziw2DldHV22K9FSSnyqb0BUoc0BIp4ENJLfQbt7903cumR5ZhOilDx6
riMtbzf3wlzbgFmAqw7xXMA0l2mhidmaYRdKKJgIide9hrVKBnXtlzx9TmCoi9QCNDdjzbYu4nJ7
f6q3JVq+GaBgrJu20UzL05vtto02dY6SPf4ULzodAftwNUiold2syhlkAuebqYI+yqaLGlLtXGTe
xmu4CQJOaMXBRTlIlrCnXQYcuApkfOAbnIQADoql17JNKLEnW+poaeHFSnulKfSuNZP5qXLyaUb4
g3lgnU0VVb+7u+qLo9sCl85+U3F99AF2gx2qdM42xT9Z00h5YQ5wo5ZHtjX0U+u9lctd7KJCwPUQ
tae7U7hajgtxckrR/hThKkaqpR1JlvmBVRgDNhEAwBFhq510JfUJpFjBREsczFH3gwIK+gLIS5fD
yEAu6hU14jvTpC22q0HkLMwFJZJnR/Qk5TZyUvVP7GAr+pe8K06UnSf6Ublk6Lsvb94QLxMJpJ/p
qak1s5EDC+ji7fsZPHDNLVBTcENQhhbMGioGvUNZM0KLWMYam5pOrK5ulqLw9k4G6YPvNLRlQd8r
K/ZXsMTVz+zXszWhVSWmBIzcx/V4owzqBrJPnlP3j2UTj4ghAjB1+DSqkggc9gyqWv1LQl6LBqMa
1grp9qXf9q28UQBrn3HbcDr2tCTgwoVb6/6Nh5YA4W7eD0r+UYHBnS0v7E1vMUb1bfsPVfJarhIB
X+ZBLmwsebJxEvxUWrTCib6mZuGDNg6tZNph3QZDh6mM9LAUg+AcvjRcEMtiADN4fPCDK0jnH2DT
03JO8uTkNhEhEXbB7ygx3F2zGzrcJ7Ltbsv2wYquqlBIMgZfJRWXw7IE3C25+KHXNm9Ut1vOOCcR
JhZznpjNEkxJ+sVKfRw6YsmoNeFFpCK0b/xtZJfI+STlGJOeQ9pyK8iAMbZHi9yqkuJ0D67ln9Hm
LVY+4FKQ2i63CB87n2Zj9HwFWjTfeHKfJpuizs1pquPlzfWGKbLGtUJ0sM0hkbWOAdwJByr7iWdR
ebdJzm7iKY6M0Uzc53nO+6u0Nc/y3+gVi1VIjDXJWu/N/WkbO50wM8yQNrFhLxNzyabKqa1pjsjY
zV9AI3s7zDGy9C5fR7T/Ga2Qz+78SXnfc9GME64wKGhR0rhrNKozNnuVuQHX40StJjBwQ6qhIWFi
U+RZhp0Z3si9b5vjG7yquCSSuuiYr1KnThsZF72EbkM9DhJvoCx1uiqZ00tqgP2VZ3nVbhJKQUOh
JutxM7vH9IX5LXEZT10YEeEUHEwvGC349KC78otNa3Kmcvlos4aeIoRHlJqL0V9ewTaHkganJW+l
vBxshw+lKz/Q4bolYXAxVLKKxoapiv6VVZQ87bWEYgYOcFXDvCdfVM/ZzE4iL3RkA4UsZvFfjdTZ
dhlXoW43rGCkgyWeOMkgIZlkxsaTpkRTGW+h4j3fZKnfQYfWi1u4KsDkuiDxUmo3pnF9Ct6S+1Nv
kOpdqE9cXD3yk0e4eGR8VLA5RFHRlK0MggFGkWgbd98+8YrEmMWnKdP193KygoLwo9LorI+Kys+1
h7BilyFVYlWvh1vJ7HJzFWbMQ1qTJPTCywVBHDmykHYyZdQibYtnENLxm/xXYfRJ425twdnHqlrq
qTAhaIVpLh/GihO16+kfMMe00ShqEk09ofDLVHr2/AXD7ze79vNFdnkHoxgE9kcQKJ9KaA9/J4qH
n+I9WmDdMHjR0aue/tzltZNiEK5L3go9ng94IkPD/CXw8zlwLB1gTpTbNeYYKVdfhz5PnatpGOeR
8hTCUNSm5q+u/XdcMmAHr4IXyY+y8wM/mmBL9XSCnX36Aes+t7tbGNhANgPj5SqdwU/EgSA5fqiT
9XfQVXaO87+NI9RUFAe0fA+zmuBLaDt6N3rGmpY4eOtrKP1esmA/Mg3kK/z0h97PkOQjBSIVBnIA
LfEXIZiYCBSl4VP+wd4RjpKdR/bWX/Sh+dZpAEZCLrwrEyk6OP1K7UfIFXlMz97GCC7AWgv6zf/e
sbCbTGCQ+wBsG0vOZdD48NiJMTq7uExVVv1XclItitXrEQ5Bx8RRRyhmn7nKmk2PVyXqJmtP4ULw
Yfy41LU+dJkzlC+H3CHf+KgE9CPQkAvwrfXRwXUCAinL528d2YhXc/THv5cXOgcxO41gIP2ufpjP
5r35l3B6bqJ1KPyXq7nHkUiAuhUQqMrGP0yHgx7N20GleleTPoIVNzjurA43Bf4GI44k+NkQOIhq
I74B+xwqoq+wKXAU6VxiwSS3XhrP50fJjqVc/3mhw7Gmb4Tct//soBBn7kqpaMkcLTcDMqfY5UZv
4vNRlyHQpp7lycHVw3aEl0BOMWMmflHx44KLd9We0GiOSuHRsfFZa4uqCaSnd3Te3Yd0wJ6D2Jv+
2msqXIPdt5mIySUedZe+7qyqSAnKDqxaqCSxIlgi9JcUiYSwHDPO2ZfZHrgsBGoGMkLyb24jO8PL
QKU8XVYrxy1IKLqVW/a6ejQuxSmVLRL9jYJQbsx+Riw7xyrRfcb6ZK3D5MmsRR8byKjJk/Z68XqG
PAIOAyZXv55VcyvYnssnwl09X13nPFt4yPTroNv08Sbo8hP+fyfuqMtzph3W7Bx+LJwpnrz2nI5j
x+m19qAXsLh3VVxFZylT2TsuHAwTd6yeJrXMtz58nRDEaXuy3ZUCwE/j48zSM9ur6oh5Caoe795i
aH3PJ0MElF5LvAJjq6OatrnoYv67+5wv6GXl9mi1KeXTR096wWPLrok9QJ4Xav989oBP77wLcVIH
qdCeNRH+Iq3RS5/iZACH0zVaCa2CAXf2G8sFPLmmdy8wISyklSdwGiuH4/pv/2CPZYKHil4nNFsz
3oK7ll1CIwFYlhSV9ixvzeZr6fhn3l+3iDZXHrEPN5RF0d2xx0x8DgSeifEUpXUHNs/viguE/tuk
YeCjFW3A+2pvH5k4bI0ZunSs9MJZK+TJe0lobD3vfE+XBN9yJ/ycKFw+3/IxGR8pIRXxARxsra7U
dwrWzqgYmxwViNKWx+H3CP18I2/dgM7N1izbOw7P0oGmrdHfrhhsHp1KCE+YxxYhj3e0reybEXOc
OQYfzZG4T96pHYulYXZsO5exot4ZA3v4dNLLDaEURc/I/HP/9I1JzU/6P3V+ycAONNQphNetbAVW
j+TT8pFpGZR9wc5y5m2E+8CTkIvFw0FSYOaVpdBT6pRqc5sxFz35R1Cm4bOJFbOABhgijK6b65Ql
adBz2Pjyx23bERKUua1aql2SgnVCIvkC2L7YzZYQnBpb1MR1IR1hTdW/gUKMzpz5IZBblhM1prbx
v+CEgCdqN/MGCMqTsOLOT69lZHcTRqggk2d7quC0pSPJD4OrvxQMJe9+DOIi5+y1OfDWyTDJbNBH
jkBEa0UIYm2smU5ZujW2gP+RZudWIXRupcLLAh39gJpcVbqy+5P5ASZLtRmh0gX1H6+rGjXhZ/5/
dOdCZ5iA88q6bbhYYoIGWNGyzYlDQeMcTrUlRP9JqVd/YgHOxJ17REVKw2/qm8tluR691M+eNLGf
yipkE4HlOtyFMO6cHsO3pW1zHIG72mRzMlbVSFJHyneWTXRTqggR6xq7fDZoQyJZkHEAFOZF62Ew
1AavTCSuCYVv6rSHI9AtMCjym8+9Hftp3Ll8JwCByn54LQQsSwbWKW+5WkH87KeLoKibsTY1jma8
h3wi1xheStaeWh35Uxfzu1gQCL1B2mI9UbYKpYuf/io0R9a8o7HLW9khuuxBu6XC/y91c9hvsdli
7LvSasrSIFbjSPWXUEj1D6fBcfuKMbRqkgebAXg3rb06g/Wr/Mw1pgXLAA2gj+J1JMlXoeGFjzPz
3WAjc5roJblNUQng5ovdbPu9fpeAYStON+IvLYvl0ndWcfWFrSmb0/P3ZsASbjjUTXFsQgSAP9PM
7TSZIoRzLg7m0n9VryJFRfiVmxv/p9EbafsZVgcaRKE3XbwK4CSVapeyYrjLxzeuy/W5ORSxq4kC
QgtgV3qFoPm72Abdh+s1On078AERE2zXyeOrk0yRN2/Hn/CSFkc+XKvqNn4umJQ6sUmBTvX4xJ0l
nj+8HKE2rKBtfGdY+xox2P6DZUCCFWe3Uul2oZSj+ctGqf5Zu7lpVAS/bb44plyLvCdBmZANPHfK
wQ1EpNgaL5SATzhZfwJjS2mztrpfD3m2Oc023T8qN++ooJAnW7aylS8WHs8S73z+4VWRq0XlWFRk
3wPDw4FRzkMtIEf5p8vj84PxrbUVAjxoFvbOnaX21YPxbkpUyPjNzv6iVDIwDAOlQbUnkCBYcWpJ
IoQcArxbiPyMOItsr0loeldQGH/9+3Yqpo7z6/fch+n/9jjDB213vlwe/QxdtKujbcbXTQ26u7LB
mCZvU3ASeJkRztgSlpbC045qphQF220rdcye+FMVdmg6VLioebPvdkop13c3eMaQoL7vS1KnybxO
bCfH5nM3gG8Zo2hbOqU3GqZKnCm4//SddR0vnhrHuMZjNfHCb5sEJIgsVwanbGuODB7guzbvfHYh
iN8XcJckz+OPN2VmG9yZGspejgkruwpU+oky5ZeBdgi+FjWczKnK28WpGCQE/kdxgUzcpfmd3lfc
dlzpazkHo2+B3xqAq3EToT52rGOSkw7Ol98YSQXJm0AjsG/g5jfUE2JuKj4fn2HTEq4sYMCdZviB
olQNM0OWgxEqPlTz55l3QNr6wILOJPzIhzCfNmM1Hru++O5+JtpKgtGe4/qN6j4iEjlinmTlqsbM
xqTCtYUuAX2shY7/m/HVgpQ4uQN7XMLe3p/ggmSeC9R4t0hiHWR0B1i+0G9pVvijx5RLyM7eN00D
Ie/qa/QrIDFJofbsn16nkcULdFbF96Rn80v8ocE0uxlQ6jquVSyxPLOHQJ/3zLs6jxAxTClz+s0E
eHr0BPI42W1/0K1z90NyvIGCCKisU12eApspqKDKm5LfpHeSO8EO4fvQ16FWwSPhb46jzFVoXVI1
VbZ6RD6wucvSkHq7be2bREvaIXqAaCuWdU/uzCDckb7DvzxxILAbsKE/79zsYV4sdS9Xjok4O8/f
TyKco0oeZQPNRMWkw1Jtk0C+muO15Ul1ItI7iZNldkD+7LEu1Y/ny0I/238Fxh4w5EwtP/G7Gu+Y
db1vZcqpeHFGIx1yqXzcbQnuuuIG1UVsgHJ8bIwFzcVmnEouc/eiju/K/ONTek/SI8OLfP2kCkao
YpbZ+ta68ZcHVIy2C9ogp1Wr857IYeG4JWs0MGJ2i5oO9IznEYeIR2jg417oUob5EeGBzeUQM7Pm
MUKkdzja7Pkw6pdQr6fDz19WvKfRhPv8HEyxHk3b6OYhH/UU7S+ph26ARJrX8aTr7H0ooyVcdUrl
XpjR4fnU/jf4s4RrJ91l9SR0VJECLFOLi4q8as4pqbCr+jDEyF0I1G5p0e06NRJRV5xH8WzTExZl
enuCHKutE6XkKiw0l8jGSnr7WPmLtqy6cmm+rmhXZVBlITi7LliBSnLtviZL3uJC4JxkevpiqxKm
iehXG2m3bBN3jl5vOUcNRtnYy0PY/ukKSNthPpcCrxTSEAeNvoEyvkx98mYdRmEGojlDVepRzFun
bw/IRYFAqKQ7+KvagMBHCysrOEqwe1wc1z8QSDK1WNfET7Am0g4LpMb7AlWYez4dfU5BfK9eRHjQ
20vt+GoGF3c/afF0e82mmuNdgqZdWPzjq3/oRNFzOiZXloaRWj1K24YhA6jk6NFTrAITUssxdXWa
6GTvlY9W4IlkvBdxvDE1ylwE0f0Zz5VZcjKI88HJSJYP6NXiA7qZuU5Mrd9e+1wMGVrjogPVtbJt
IhmkRojSsfxLaefSI03Ki6txjUe7fc0SBLNL/51G4OL1kCC6PEfQTSFkYlfjc0Cmm2U/Q3dYyb1f
lKSSXLpR2Vke6fzhci1z1YQwwso+qmKS1E5mghcxs/EiNCSExyhNt1qVXYjgm6ZSGzLGXyGiPNv0
Y1Kmv5UUIcb46oW9//5ZtlBxXUHkCysaGMfKdeQefIEKIKAukvL7K/F9C+1wN2s0MulZR74ERaqa
ZtOqBFxonXcYcnPcsa9tDL811grv+oOm6u2REWZQdUiOmxsS8d0IHs+b9WGwcWCFpBMPQTBi0VYd
RunfVf3VLrt41oIpEHXzSdKLy2e0ZOclsPU9WXl6ZebBwVFQZZaoprkYveFSu/XAQdCScp7p6zNc
GvphkSy6jwDixCvO0uom5sC+F7AJ4ogI9rE0EzIYm9iJvPWekTtqENLTBxvNgcPpQ7pIwnxCku9T
KDNFVqHHtwicBwezrOhhdfywfD7aiNGtYWKJFwyXtOvNd0nd+0LfYttEyyjbSfB15CSP7aBFExoi
UNfnb6GFRKLifrFyAaROqN5ZqYsyaPuGZk+ZIFULudu4HmsjKYHkIkn62f+Ic08IH+M903PaSPrr
J/e+34qXnLAIu50wGXMnyfhWWwLjICC/kngn3szXFO1QkLDTYudq/NA8roI5JJo0WJXQoBeOwEUb
zeGvlakr9Pzz/yXsNVf0ldE1M/Ei6T6jQWjrzGfUW7/imYijYa1Y+WxrWrnvhzRUtBGG7tOmGmm1
Nspw4rm9Egs8+kQIkKRJzzknkP2D17jVVB1KUcwhJcge70ohp0Nka5enBBE2DxdIX+3jFpj/IUgt
Ln3u30TZAbuVDfpyCq/ntYZjB8F7wTxTHSEisBXtwWeqfKH4SnyJBn1JA817+cH1OoBADIofLixv
0xzwnNUebZlE4t3JuMF5Y3ez0koYjRC+lC++hSgo5/+zPBQ1BQpITeUXLRZdomjNZkpTcII50qSm
SMoLFKfckYHMlqOPSm2V81PG6V5DMq8cdDmTGdpcdKIBapWXCQIrWi7QvWlbRAMnBcRZy3iG9jNS
7l+c6LZWw128sBDxSWPBLIs77KR+4oTpr+HiE1JSDJJq2rKvav0jjgoAOs/LeD3ecjdhxQdFaZg0
TnvLEy1yMyI4YCoR4e2a7dr72AL0Fx4vhTfX2NKaHfk3TRzNxPZUBqmUmjIPyWZODNz7lr91/McF
FUexk0uMutrukqaNQjHjnbP+4OuzVmllOlq1obrP2p1GNJZu662XrhIfWwHAe/GbeCYDdUcv7T6Z
0GGRrr9omBOiUn+TlcJXsLy9hUiG9+wPiyN6bU2A90uWmnkdjDvYQ3qx0wjC2PTd0VizZsnMcqB6
V1hh3FLuE1S+a6kjjWTVUl8TvOJYJIBotCXVtt1z/hRMAEmgh2/9vLYNR8sHYSaB6ubeyLzjrY0i
PH3F9/ndBFOwQ63wbG2jR1/jNLtgw2MftPXFmQCTEH1UuykqSNhf9cyO/omP2jRwkb1gU5qnsctV
ATAkHoqrQVTRyNWCiuHEAPU7zcwygOdjgK5of/+KvfHVzFEayCICmDLXkqc0PD+YM/00+1hzVnba
WAbH7O6XUHWCL1vCvrFIJ6yiN1yUBAthmEQcmbTFiDGXFA+ONo0v7IkOVAcllULP3++gR2RvJfXB
Sp7r4CR0jjs9J6PoR1qKCXaaHzrpcIQtJ91gyK1NkXi3fTS67A1YzXWBU7ISvF9lBFd45p+UtUZj
7+o+HBjal345V2LOp+ALOKo2CNdcNQqDcoQ0xChTv6Sl3kA9wBnChJV4eCC3T1oSipKVbbx1+VaB
xOE3t/KlUUsAj6wXU8Bsn8ZgvGr1lrqWWJBkxLZtOgB9jrXpecmMYbmSX2bIIDLArdM0/sJmdVff
0XWbtTisGIGtC77Tx3FwqtolSogKTMXC+XgH77UlsYUyO0OL1CgnOxFdIgC4W9JcE7beCvUl16N2
OSwQvei0p3YFG4gj2r7HVclKKxcuZubOso8p8ACsSEpQhMzwyECbSWz4dOnKMJRenroY0EekhoU+
Qfjv+VdrUAyAF070KET1ZoeSOzFJvBM1K4sDbFfRUkTJg/+Ehfvk5TjMp1BVKUYi8KR1J06fcPeo
umSQO+pHCQXdJfCttyxx1NyzoItJ5rygytzYDxtoxZ+k4Ce9ZolgctSjwB5u+2Z4ltbdf4bSQpY/
fVXVCBJNInLl+2+Pf8Bb12A0s1f1FuEPuiDKn8vlBCm1vF2a107DK9LmL4hLxxcBrAcqE78aXwxm
e05bnyFJ98GxoO7uCA+c0WRVEdEFnYduVtd/0xh4Vjvj3PVltq3yAZmBaxdVClYerov9vrkkAMil
PgPnG70vtmyeKmDZB69zzw77bvFHaFJLmp5csVNpe5sFWoS+FHtLz5OsyVtE2q0sNa7SggT6zv1/
Kap83HSLx0V5ff/GswTJ3ZgtOA3eBx34wffmW/CxS36wxZhRb44G579MFyj/MmlcqyzyRUHoRC7D
b87xm4NNIJ6oBi2cjKZqThG/srnbpYHt3T/bKUKIV2rByD0aO7pfP7xr6sKZegvs6lOJA0y60Kvf
UnXMehKd+p6vIHaw4/ZRS5D3ttFLNueP37UfC81Cl9duGkLi9RdRk3thwP3skbSe2cWIv+swN4RI
EnRYq931ow+VOgGOAlABRiPAtBHMhKemDEJsVIWc98DmqENSqsjlfhAjJk1irZjwp25lebW9R5wG
3GESaFLg8Mwa7LBcZ1QA6D7FjUEV5kMgy0cgaImrqkozo09hpfxe71uUwCJ1VPal1prpJcFRn5J4
1uf7VHreO0TpFg3VieZcMsV2MFqRicgA8bcqGiMbSfNd7Fq5B3DFsJdL198rFPCG0gGtUIRJBPn3
zuOSre1MG0NmYcddjYg7VRIpWjopOcJs+CJfBTrGD8/hol5LUQOVjjs2FUV8sr1bmH1wTJRMaJnM
X8EVYNCuJP4eG0jnuaDt0y9TtAtgwvrh3UbwkFHhiolQ/yGD0IuBk9GOo9zuWzSU0FrMnSLcEzG1
Cw///+043Mj/S/VxJhDcjD78+E5/yNxmbfPQ1UPuGQsF/PFHQbQV9i466Ca6gsAYBsYKEnEoOKY3
OSXaG8y8qrV1v2tj8q4UNqhJHTLS9/kxGOze3ylR91y0bmkc+e4IEoFwRuURfESTj5jDxNbG9Gnd
3feGLOVlo60ZxpmWs8lFahwypvaTIXe16Bx1XAh/JsIC/XLaomuPJecBZT1h9rANRD1ooAFW02dZ
VlMWmdVKaFZiD1BRJS/qUpYxfDf4MT/41uKE5NfhS4EKNEar+XiDB79ob6Pl0h8i7THPr9Spy2l6
fifh2shyAut8rfuTSrS3q3zJJ6w0sGcLxfVsSUiWUs1mxtZyO76vheuk688lyj8D9CX/VsQMC8dd
EHzcoxJIXB7S36xfejoHbA2ig0BLV/HLGAT6vJZKHCyYEQlX0vgDVOO6h052DUarB76cQjtyU+9d
s/bWvfiSaMr+mCBsQoHYkERZkPYrgIVJ/qR+eEPOO9vP0bdHHC5y60qvddQjjtigYsWoQk+R51ib
cmVRJWDPnN/huOrzcX7f7eZZ2xQxBokJFnAiP0WjiXaBV900yFAJ3V+x+8aTK/2DSBSv83KnPCvo
LrfULmzcBW8zABANKWoJk7rjnsCZpoPUCy26k0ynPsztr2q8Z76cgWTpnExk8vVKfWt93jre9biw
F603W6g68opT6mKQqn86aIJ232pjdBlt04g+OSN682rg8XSRlN3+YmI4t7jQnb7Utjvk6uluKcY2
3KcKBjrX3ONcJyJtBu6wK7ORhzndKNEc3nn4yTAeZPHAAVySj8rjU2xs3CfL0LLr54REAldYbLqx
/xK3hxTTz8LusJXD9WQ+8WL19HTmw0zV3SjczkZyGNLTvEBdlIdZsUoFwtErA+RjIP5GA+45m7h8
CXuUhku4JWW4GDfWqTT219Ikols2Ux1oNRMoY3Z/AgcFyjbeSlpR5sj0bmgooILK/ymZnGJLvpaF
2NJTacb+oMl6PFxY8qDm5q2GKwO7jdQ7lBnxtmN3SCMPChoPw7xuxyoYuYNuYEmPPvB3xHmOTvho
CuoqWR4HFn9QOEvipgNFJcjPrHZ4DuX2gnQpECzTM2XVWRBT8EKRS3ONmuDH6yM7FVMWuth7PDYm
Kq+T+tRZb59XWlroJUVRcB3ocBN0Eg3uIm4qn0jUHrJ1C6Nx2d6XGSBRhI/A2f+T0niNKC6qXvOg
MTCc7UBNSmHDRMOfx4GfPlOOchOYH+DayFb0eOmLnt1YJ/ZHzoI4JBuJ5/Ms+8MXlD0JTF8IJQ9l
srTsQRW1RdgCafrGrCosR3AIPSd0Ldw0O9VXx3iEntKe6gwVXGQ2u3cQ2bGZbIL91Z3hQGhJFX0K
mwCIG5qWMgSSS3xyCIelXYSujt+dKINH7/V7ErtnKaAbfNEVN2J4TumyrrZT6LopAzBX0q7RrN91
m8ms2ya3XeT7nxMz31tI3512NoI33En4s0VHCqdV2s2HyqPRH/sehVvF8BClR/yUDJrxFbWrOxJ+
r/7LiC1D4sQTbXYO+q/xSwIbsOIrj0/pFCvSmUTa/D3tk786fjcl2AojMMW7W0DArdes6+lHQNfi
c2idc7qlxeSUio41OCaIQsX8l7yXzcL2HflcJ6pZG8H8ojPZSdrIhczturdbKs8E7RVqzABQkKj/
KYbdw1gmsUoluf90T6b7CClIvJ0d7QhSDRxHK9+44fnI2Byut/Ca+Eqxn5ozeTM7I0vbjKWqPJca
Zo2eGYxgsEzCav2rXZMoZm6Vs9sEEOHQYQvboCRVDk0X+kSW4hOYWQ4fq018yet2+W9qvt5yvefs
WBO8m9ojMspm7fxdAmIIG7wWUpRNxWSUxiPtMC75DbXs1hV+dQkN51aH4AomvwBb0L7biU5z5hTf
NRfGAwcL4X7gPAFIrQdMlL7I5Lmi2y88TDrEUQaaC9wr+yY36PKiRHlWt7aju+lucmqexdtJ15UH
siEBuKluxQYj8q5KGDhXcrDHq/MBC+p80gUF6FqgnFEvg0g6Wz+tydQRlmlXKCPGhaiK/GI+ITax
+/NQeCP0n3mmdT5ZiYGwz/X+poRyHUmD4Br7AlVxpcp3tF5fFIN5EEWwhKVV+UHi92c1if4355pM
PNTgq/+EAw8FUIBp4YNezuPpoVddtq83WTd7LU1b59EZax8JFV/K/HQxzhHDRS09z+7O1zKF1Iox
op11i82qhtpBplt3aT60a5EPPxSYzLh98secxFZIxWOtqpZ/JEdE/rwcq2EoUOzWUq5TW5QoTdgM
IledyrgTAEvWdGiQ1Cyy8TKXr+Qu0M6ibGsCtzwFFgj69fBLIPvb1215EJfPN0KTWXKgAzGcVxiK
KRFOfABE3nBVtdHO6tCkYSKPGu/PNHTfDK6gx3TtbwnbGxN9OpBaOMMlBE2hm+IrGL9tlrcLh09u
fCgRV7acWeuVj0KzEXlg0d4LAZyn/dFLHR1QWkVtdGbneDFb9TdWxZnmuchIjh6X1bxwosH3iiZK
XyRdt9U13BtMnc7avSgRoCvnJBZN8rCgN7SH+K6xPj71beX54ewgGX2B1lluXpSLRSPisKX1uaK4
+3a3+1mmQkVr6wZN92mfokojHLFkY3xDWOL1455S+YW8NHdXfyLPHz07a6wRtotPACa2yDpUs1b3
s6KeldW8WKqYqbvOde0bRt8wx3NPM+vZXnsDAGos31JO8Z5abLM9AWmkCGJwZhxeoQYRElxjXsid
OXCzCdUquat/mulWOHvHIZepNtIPcN5iFrMazfjqpo4T9rCbczbMnJrYcjjU7S9ZQkUPm3F0GDoi
m3RcdlM+jp4K2debMtB6wT05Fhhz8Noykew0R0rlOooBUv7xAI3qdQxYgWGaaMgsvgXeGYOkClDX
QHUmwjkGl2cA1ciRGaPuI+muzekEMRLp+vWFSCjG2UZ31haUZRETD8jPgsqunALUS+A/v5DInQEd
UMAOnEeE0zl2t/IUWWxZqedLjlUqbv9mJPOOofcttlk+nQiZqVShMUF/dEuI0Q2Eh8+qbmh/SSsv
RHy3kf//3MyQgaatbQmQtm559sa8TQbOTWwQbeEb6cqPluSN8Jge2XlzTrN8HNP+IVkeayQOwzSi
dVWROwtHzGsCqsFTGxMU+rk4LK9TPp2BVKxocOY8cfk+eKoRCbC2ghO7P9l5a3MQJvtpWCZWD7Wv
bt9GM2P4cj2f+tDeU9BuFQgVZfnXPd9+kGg53t/24/WAPnmphx0pF+NAZ3ymUvX26U+TFPuXVH0Z
7vsvSSNcWnKeWix0nnOfMZ7ESHY1is8sW2hEopLjVwnPicSGS1G+ekQmkZFPFYvnyjNSTb6E3CQK
Aui6bE2ZUZT+HMFSIHvGYrgtOSBsnXv8y1EPh4cOeOR1kwWMZZB2zchKLAL8xC9Wj9ux5slpj7FY
TdvnwCaZ+C0umcjWflq6Kep96gZmWdGoPkUwT8qYmJYaX8GvAGoBJ6yg9tC/7yd2U7ca4fkteSEj
mF24deAQOx6kqvCpfD8tX4W8SYrzGdJOrBqVRBLnLtJBI1gvbB+lZB6MqcOoyc3lJ2b409kShZ0Z
Lnm2yWz7WYyCk8IyKzNoRQqejRYinsum4gyBwttD4DK48lPvLugFqNQCJJY6pVk7eWu8795gzLY5
9PoVtDRN4UZz1+4uQaa5ICy36vlX6OZduq07GF7FbQuE0eZSEFjwrPTZvbIjTEBsYqmZmqtiiuSF
qoRysON+OyhVK1Yr+Q2lOrBS18DcPI0IEUseaGrMoe9M6cDJ10q74k1W1SAVmtr5m29OLgfeZGFL
zF+gZWb+NNxeOg8g/TqmPBwExGeYQR4Ru2vHLLbYYyfK8tSRheV5NIppBUnuZnkVl1pI6cLeE5mD
qlFA7fQJ28HMfdVrKQtiXyj5Cp9VkfEQkYiTuutGJp9c9EfdV9hF6qmrdnOL/sUstObmEH9lyJzZ
AHqO/CEvdrAkTIdA4yn4gva27pZqyeEqznpyZii/dqCOlkkzPLmmAYkS4+lA43Pfajga/j+RuLW1
7g7hoMcgLYBetXz7lljMV9wQ8rCT/tbq6c07Sf8ZSZG3e8nqsG2RdALpb9cdQgdMP9uFP3qdY5qg
oboiFdMjP6rwE0kDjVk04GycSs7/bl+3uXtBvdD/6qqmRXRn+Va1iFhUNo7m04J6NzPhxP95E3xB
loNoYa0Mxutbe3FPFF+IK8Jm5Zt/73HQHqGYtUfVQmKDISsFHI4UoK7jVJZIG4fun1uQw0Ngj+ky
HsGlaqLK2AcXVjBCVElYex4VonpOXsJrcVmRMnYoZn2sRnPvL88DbAY+70f0NgF/59CdQqnb9jLJ
geDx3W5y6ScBya1DczobO72nECiaWQbA+ugHbgsrdKdGvdHXMUiUuTumZGXSLjL0K49Orn7I332Y
a4xEflnU2uE/De3hhd+xwydduubBLLo1lHFQ1PNjzlAskphlVsumVoIhA3cS6mCE4d0rdQwq1xE+
ctlmGaTzKs46kiDYvsnw3ToHFbd/kvy1tyspIFP0ODNo1/6mGJgYnswwyRi5gFITrjfd/N2K/Op7
w7/ec55WDqm8f5zEHVcvWZdM2EXSBrGWEa5C40MIWndalAZyhgMjteug5BuimWrvBf8dBcAuWn7U
2vprlCHTVQKdMIWwUmvb78bd6FzMk5rcsi1kd39RrgLUzJYnDeIeUWSdcSO7YoyPGxc3pwYajy/c
/FAgF5jMWUMILz9Z4Ivy96aZ+/7m0OYTjPcV6WV2OiqFWt80qBbvQAVh7poRiveRM7KCgbK18EHq
8AovOZVidD0X9YWyKaRaEO5bn9LfUCHK/So5JHDB42utGxcgyzbK+us0sXr5q3NVtk1HZRyTjUwG
84qfG2vAhuUrXyY7edIti0UaLZAJiD0SG99SSSvcPEvWB19kM8Q0YJskZ0MCvHjm79KnDkqtP7SK
D6I73yHjt6pQA1ismaApJWGKGL/6n8sBHnh6sASuY9cKtoYtj1QcVO3VLJ9JTFnNGqNG72MUVFta
Hf6mjbZZptG0zqS+jpM0INpQNB2P+A324hyoWugz6FYlPa0MffTYYIeo9hyVWKx6okoTT8eHaRJA
N7bK/ZoqBUoQP0WgiVO2rjNOeIR5YW6jofOUp42RqI1r+YugmrdesCHktYNet/HJ5xuaHg8JWmWn
dSYb+JiPR0KmQOLP37hKfBCA3/xKPB5R2+Z7g07GIRwp130+PZ/GBrn9b8gemP8M3TsI/MaBACIc
OQuEdb8899TGL9vEb1H1V3J05Y+2r8gsShZaQUWL3gyFe5qVgt4H+pFSA3leO6JPwpIUPVdTy9gm
ja1y0fSGK3GZm4oiAsxvZ7itoRcfF6xrNfUuIADmVZMeu2SDLbGLwKKN9vp9WPeSVi7rM5r4/FOk
SLJg2mrokQT0TcSs5gE6ozjv1VQx/psQwWdMoC5OVYP16lS+LjhywV1qMUQKIESQnDHp8ZHvvYOX
F4pCxJu9d4m/t2/EIApiLG18Wg1oRr0YJzf8441oRu+CB8Yv4J4F0oyY+WHdv9yMw4MgNkrehI/X
jIx/j1gl7/45dVQjsQSf9gvCCmQxllm9eBYVU5lHrXmnocncANQeDhSRgts82308BHvYK7XhTP7e
JlPpdyjcJO/K4m3kcjOKVktwTAWlnmuCROPIqG+9DQ0+qSWMpkbuyXo8zonsxB7VDrT8dBOBkr7m
nw+d9SNPQtA+2RVae/SFmVT4FL69T1ozDCXzA41elagB5rH4ruqN0XGt2TFTy2g/S8TzQY9Th2/y
knl10Yj3Sf7whxEdRNOh3ZN9eH2poYWp1ZVuCHb2XUakuIlgvZRsDwqggmeZnbDYx/ZMGpWmWZ2f
IgH8qASFLp6X8aj0CCL/KvVWYzH1ZmgA9T0eJmIb9WcMuEwyRg96h+/vlcr9/MPmkupYVsUj7kv3
piBhtvq3HnUKnv9ivvdorwa8NgUEnyD2gEbD3K8tko2LH/1dRdccO6q3Z21EDXi19FQZMZ8i98Ee
O4cUTuklNRU+JsD2u+jdaz8UAIVscy2hO2nvWdnpF5yH+5Ize0msYzysXnjO/EYmHgW4FE0t+8OV
XmIBPpLF3Nx7ErvlOrD0mgYsf9Qplq9stYcOKYOFMesLSshNhpa5/Ao3QWNdA5EKuRCLR9trLWrV
wkl9p+D91IuG57iNVsK+Uz3beWmy/JwDbZ+ZcAMWHEGwgyKaxnfKKB5Yd+3K5OBY+kaYyv7yat5m
wM9+lkAqpe+LVv3hOLGWph/uMtsublpRyU6+fpYc6PgwlnEVV7Uoiu7BaC+ZTia6epxXipRWBaAW
IYrtWq7ze8gKZs+BvXnRAXVffWeC7wAgv/5asxXg2ApZ4yCxSNBBt5IA1CPDomcHaPk8jMWqXTQ9
RrUwoqrtP1bC2TaJI4WB2zlFHmueLO8Qp1sdLh4r6m4emdPnlzwFflNt6ZNzXstbm0u1vUzA2gaY
l7+urGuBg4ZaR4HzMsT7YOPlKPJ/cgu7HZeTveVSRnbyWl8hTh89v9EFPXza/CAuHTKoavy/DG1A
8KnibqNTVDEYO7ZstBmPuYoiEWdlTatdXqlKB4pu52EPM2WNF6jAiSfG7Y8ESLDNuqiKQX3bxxnT
SYcLeoWwzl52juH0buudtPYx0DQU3jUYPNBGMr7UvrGPFWagRJPJ8f+pqfWuG5z0JzlZVmiqnbZS
rGqOJAHGHgRVSyuGQkZ7FdsWtBVm6Ep93u3AkBVPQvoQqHsdkWUGP9nw5wQN5pYBTk12lKajzKVd
uEn6SW5/ckuZTgqQDIuiIocyM4doNScBOpyHJYP0Rci7JjNXZcthLQMtzHCeD5VqoymjXf8O3w3L
+PqyHo5OMJbyuDnkegonTLjgADZpcfYy7BFI11qYZyp1cz+6WBSXbv7DV+1xI0sl1GsPXapvdpwf
//4qNlGCJDMtuGtggJo3H4+OeKOLaHjJy3b10CnW2JoWeJsh22N0U83f9RYFvVwHgeyYIDl0E1lf
W1HjedsLcp0+8xNyswA15CuRhEvuCqFkUl4pbGnr9JzT1dYO/fQE3HjQ4LWlMLCNvtdxcYJFVbxS
Z/Tdd+dFpsqC36yKbrxCOjeJTlCCcVIJ+R7zGXiJ56MBJmQl+dkEfJgq8hNXpRfvxu2iBnyR2CGb
5L6H2IoPpcBNUDyl8wmnGiPpnn8xTAq4JuUzPuW3XGUz5PH6BxIPhE0NVti91uyhg7a8XJEdVief
qOQr+o0sHatFt+xoRUWlQNEeTn2rbarIRFeQF9iDaK5f47EYvnf90pQAMey/ljyv1/c+goFueqX/
WEfb3X6dnltjm915mO5HP8ze7zLPdy1YSfYtrBbuR+S9T8I/LVaIY+390ARFAEq+dFa4quDqWtvc
d4+oCBYNscUU2jhxtPeVNwkEVJm3kL5Evyeg+GvFBE78fnokCqWKz29J5TnySDRkeqG9cr1iHsI1
Md62VXcZQGoGL+H6OijeO89CPAXuTDefnd9ol45A3rNwii9jaFDqfh211HLqIhKTWgCvXVDUDOz5
Dhz5IrLbKjruJ5+wYQmNJ+WdQhau8WHddq3+GDX0po/oYP3xlMOaWTOoupgft2kGP5wiVLSenKp9
mLvb7S5kGGOqDzgya6x97thuzIJxbGHncrq4x6W65i3s/I51MZWLOmxh68q9tMIcE/CmufVuASeb
qUZ+JEP8qtzcsNR7/rtyiNHAPWPnAoSn9TmvVxZeNs0QlZ4eS5upJTVX6/EiOpNsg/yJDbV7g5DO
PkHQR9Wq2/odChyhVy+9eqeFP4icRAHvv6lGaGczuvnQZzYfXgQnr7868rFPkTMaaREkXWzYhXxH
Sv0m3UBiiW6sKjsdVgtcz0N01GHOuLqL3UkeAPiENiOEgqKd3WiUfTSURtO8bNBIko2G2xK1hMqQ
AmQCf/Gk8+XlKU31aXfQlTcnCYl6UBeOnVuq7tUhpr9vH7nQDe/UktlhGUyUuGdVac9CXP933OwK
tulKNJvGvaaqbgYo68yaZqTQhJkYjLn+frGSsMee72VlyP38p9bSidBfCrv+PJKTgsnlGHZPfaot
6hmEywuH+9JM66m+FIp6bBVxPHqGePJeqzMGhEbOeMHCaFq62nruQkP0qu0khHj4kklSKaz5EuSs
scjNVE8xPagGBJnQJU35mUCLeJGePprtn5N4ht8CqmjW8qscAkDlZpUOHZ9aWn/T8n8or780ycqk
jBSfweZHJpMeoNyXqZhsXENcr8a+UvRXtu57ChVtVSRGbJBAWYMVv1cO+y6tsEn5wMgHOxBlHmHm
cvIOoBLrAdHndmnHA0Z42VOlxvlnRQBwHiX5M+auZ+vAuqp80WvbzR1h3t0TxLypSz5mWb+mdPRI
+i8onY2nIgYPEcXqcbpaCRdUkKG1sJNvN8omfc7HundK9XyYBXHigYMILaWKyCzvtsmL6+Yi22O9
cx1wYiNwmi3z/OZKxqR37iyQeWsddWMLNzTkUfhShRJAjqRcsXNVkYTVu1lYdcr7Qb+BFxnS5Ngn
jdzh+AWv7ihH+xT09ra+4tWKBXfkV+5vh67knloYtWQUUo+9WABVz1qoap+p8HxxwUjyvNkebeu8
g0MFqqdoqCTOtEhuo2v2HGQrMWvsoNAR1t7Urd/nB5MLOnm9wgGWit7HSHIA/s+qm7nS94gI3flr
V3eMh+6kiZspgU/WN16454SgkGZG1I9ybCgLi75aDIIVITuOCI74GGXl2asIsC0ZGyna1I6ijD3R
Ne1G5+W27F+gm1jcvycdN+ctQr/FeyKU/rDeRIcIDmbTd34q86FunY6kWu6Yv0hLpwiXnFjKMUaG
oKqDQci41Bg+sy8NB6JIAfIwej6P/0ivJsl1t+ZCA45r2izkyt0MkQ45B/1pDMkPKfAer53glLcf
ll1BRBwG/Rx94AhhZ3iA5aWxR586XGMoTIrKDbiAzmP7b9LwwthIXxbcIEncLWsKVN/Fcwou0psb
D3vbVTxDTOgm84nTQFDrRXA3KPOb6FpYp3cMrpYr85H0Xi0ZR6GFcX2JXT9m9SglZBcPwq+BDNnA
nwteP9x128uWe6j44sZNLGRQDXrG2C4lJuPen8RpkGEgVgC677SqQxXKQpe5kTtVLYsbSSV1K+bx
YgCpLOm3YPoAuTbMkMzvjr9IRlhlglv0pFVY4vX0uuPSMIX59AAE9xHJ2s506AD2RhD7Cr3VRb/s
1kcqkCPCPv8B7KO3YsJzIpcAU8glmA/7HYUiQv2TAhgSyddO7fY/Zoe+94W7XGEM5Ef4lXZboQK2
i5sG9JsI6F54psiTEtHscT1boksU44dqgFbXpagKRtD+jIXkRVJGwPZHPLiQlb3R0stEl8uEcYQB
cwWwul5+7qmJz6wfuPRda9ZGE39Vpv97w/y21ikBc4PnjG8Lfr+wHVhVSV0T3LcXnlk6SXROg3i/
GiOsTguIW7H9DAXaeugrcjfYRjD0IXjx+/jFBei1bUF5gGYxa1j9enDG6txKtb2yRTuNcWd2Hszh
iRQGHPuKO+a15MAeNP7wSrXeaFYthdo/14B9lbpK3DvENd3JTrRUl73c4ZuZogsuKNvx7o9tusdv
kuc/f4PAe+MQzHpkmLV+M97M342O2+d/62FILy+3iIczdQ4enW38WI/H4erPyvGb6sWwEQQkV6L/
uTWYMJiZyU+192djkl52kji8GFWD30erh1W3CXzpwRdkv9mZekM4eOLBgZKOdP42TYf71FBSYUKh
dwb12qOpgCrIgLG5JoriwzSs7gxnzCUrfyv9hWJ+P0uoWcZ8uQow8MFKnINgHe27hb05NbG/KLse
/HWqbfpkZF1PLpbjtOlXgmelfwnrcQNbvTa+gwgc1wL+W8iuH2czpPBnjsudk99yi+HdUKtbqpsM
0rHeGfNkRRQhNvK/PO0ztlmpQRTWnpkNhCOru7H9RHHENJ/ARu27Pn9oWV22I//JXU4D+Ck9KezV
648kbPISnqfr5F6BbBtD25SKRGrrFo3aCaz0+4lgAD6Rdsmmf76OAmR9rHthT5erH7aOlh8G5hP6
xakN9T52jIRb1UT7nlFcN2HqpyU+Oz/ym6ZUjFkzrPYXMH+fXclC9c3kSQi9DJHrt9dnKrYw7LTt
tO+woJ8SENA06KOTNU0eLJEm+Ri8nMqIhTrUIfFPXsl8X6k1TyaEyqFAqTQIQ1bg1O8CyCEeyvKh
/NBjU46J0AOH7yqzOavVizqx7+rAXAL7sPw7CoI3c1EQm456HBJnxcUalhobZuo1qZEUW+I7JWtx
IzcUZzcrYW4rxWE0TxuU91Yvtex98Nl/BQnOjZaFCobMYs5uLR61fCJLmwMVqaUFRVKwDIVye2gP
q43oTz5fy5cDvWyVeT9qvKbW7if2vnIS+wmaYH5EQRTftyx4I8HlU4aqwEDfrjfK3G2gsrvssf8I
1hxXEjIP72H67jy5hfcoc1z7o+5hoHjaoPPUa3SSsn+GoZBYmHu3E7F7FeZkuEZaw5IMQHhNt23y
1T/DEu6aGSigh0u/yZUO9G6fvkq4QkTE/i8fwQLwgfwAyhDlekln0WbFyIb8nQwJysu80I6azguh
xIh8x3/ZI93+k5wLuuozkmBOtABZv8FxWypLAKnz95gsXME680sydUAud9AwHkstdWgOD+ihPx81
JZ/xaNtV2W26fBr48A0OWUsva5ej5RFT0kKieul/AxwPaaGyu10uR1PUdPJG2/I/fTKMjqEDk/cU
mZXrE2A6k+7b0AojqJCJUReVduZIVf5s38QuKTnoWtQmJ5TkmlXTEyHifPk2sOL0ELa0LxbOQcRV
8bl0+ePnqTAVNpmoEaUqR/j9978jW5VJ8tufy12wValWAEnb3FZ7y6Q6sVH00yo1sYxAZQsha9VG
C1jdQmCTbjR/VHTwtxgYF0pxDlgJ066RNxPpxx62cCywHA9xhgbyFUbxTRfyQHTP3FqYO+zWCVha
HyyCyuUX4oIiBeCXeGYjqVOLAKoVUxglQiMojSpEARpelmTju4df0pxW/MiEAXWcibJ5w2izEGwC
l+u8dvwCIxYn2lqUxUYEugFQIslf49gHf/dFOz2vxMsu0usSJPYrpVPG+03OKGYl/vIKEzW6ixPz
i1WhM4o8MK33JExpbb2EC8oleoFh5o1VUXRIzBd0u/kX8+x47/eutjlPOeukzVh80cGLl1Ab/SX7
o/sc9o4u8Aq2EVXEso2OGFJs5vE4oWeZJGWG7UDwz82UCyag1JCDWojwfjq8lkmr1O9isQCoC2Ci
ouLFuMOisZ19dnDJmod2Y+VXw6+ym26gSrBChCrPgo2NoFujwh293YfiCdOtx4PvW6DZyLJirccm
XzUoXwYefiS39p6zadfdHKBasM8KTPCaWdKYABlgrnVqqC7/X8ZD5hbdDYZHjdkfesLKc1cwdg3j
pyjbxQ5m8yMEwqssb8beFrtl9ZwvpqO41yuIUnuwtV2Z5KXBy83ZtW2VGi7DPse7x5K0UxAiWVfy
EMu9I6RfldAnPnpO9ylcIsOlaEL0OU3D2nSflBZoe5WKDQYnDN2lPyZ0aF50VZRqdjy1qk+7Dsig
6kS1nG2o5zwzd3YCC6XOYyyzl2S8hKum/Vr8qB+UbYXcC8um8FJHdsRFSa7SHZus+hmOEcPo/khy
0HzgQ8TxPGoVb79LVzN9xMdYl0W8gsyWxfEY/Xb10fKsNsCIspu09WTV7FO64acBvU+gyHCkWBBk
B3uGmlU80yGU+EuPa8xQDJdNtJeRKNgvdRWLFlefZ3aJDRdC5hvO1Py2RdMU0u8PtYRqM08PSIKm
iK2/VHJ6hbsZefGOvZZG5jON0JnF+xcG+5r/OO3Bpx0CNa+/iuYIiDPOo5asiyaXVU/kPAXGuOF0
Sg7kALYIr+/tfW0lro8LGBx8qfk3cldM30+jmcYxxD+/Ja+DZCudbqrr4NbqK3ZGFuEie0Sorw3S
U7XubD6JOxEBmUzxYT7BbUoPvZZ+uOOHR7Au31he4lBXb4Hgk8K220WB59R9YeNRwSvIZbxgNe78
qHPXt0b9GwqOZDsd+Yk5IHn4G/2E6Zc7niTjfrOFkuhCiwzHiyphYOsXJTkSQdytpisrHiBZsvx3
La2hKp1hnex89oxTBpD9DLQGzT3ValqcZEAbyw5ytqyIUBLj5nEo2Ttuaiylzfdz3mlJjdoxxfOa
JNOY0t0A99sckFPg+yhNXRdR5jCu3pGhMZS6rQHix4urUC7kaln8nEUuag16f1KKKEdFVCZTEqv9
MbaMBLs7y+7LMU99o312vK7YLeKWvJTtXaXaZDh/mUq/+FvraaAw+l96U/hamoF4TIrIRrgdS/QJ
TT6Xa6V8N3N+t5mRhsXHY7Ic8pYYj8hDqqD13+f5fT1icjUCeuJH4aBhSW6ZdMXCr+ZZQ/VODt7z
fGX+qLJkv/QEnhxHmgRhV3e7tjb4jQpyKQDI+oA1MMxZdH8aRsVvy/lrR8fVH3H1NBaprbCOFYos
+MPSWKAWilqQeVhkbyu47uuXBqVFsN66kheQNn9NgFKJXIDKfJGPhN5+K3ll1SWVVitG4iZxCxZC
oSMeCJ8MI6CxpkrRN9t+YF/1/Vrnm73+Sz/1VwkBwH9wVIqnBDXvu+T1U5342K3W2Qm/u0WcTLfm
70Vc6VHCJN603NminkU+fgQODFOdsK/Xf7jcAJ86Rn/YeoK37wSaJkK1fnSXlQQDzZajes3KNTZG
vR+247ZQxjAEa3AAxHQm4Sua0zqkUTqHogOyBEZ6mp4mLaG9NdEJQSrk6RD6Pf/Ad88eVskjaFrO
EdR1b40oE0inUQL5srO4JJz5u0i67IpcKU21c/eASF2FcukF3q0SH1TBR67/xiaNbNmaP6Ybes8w
dNJlu28CbzeEdPYYIxr5AbRPm2bBtVAFW3IH2KekyHuqKiMgLfg3DmWc3ziyGz3m/3Vryv3vkAxY
nDukx95DjzjneOm2WxFU8UMqCFQar7iRpVeJxwadyu/n5jETpIJM0GfA/SDvmoirM+AnijcjdrbL
buyPXoNPuBlPZrjAF07yoseTay546L6a3lZ5m6QTa8R0RZ0zJmaTIx1lqCYz4ywDrzrPrICaas2K
lvqD0wkwZU8Qb4W5fEGURv6OgxZpOgr1jyvly+zIC5btRnR1osNMtrOQ9YjLCeoD5gM8N1p95iT1
5d7/JSg/Kkh/RShXtCgFa2oQM3SEpN/DslADVWXVVH85VVbikR7EP99sCsGNM7H4smnCxBIztODz
+ABDuVXqRF+fH+i79kJOzBT10IsY/qATe6V+TiXba7ZkC/NSY1N/1WEDdxQ5hS57BU/tplZUbdil
SYIlrXC8Tj2CHI4rq5glUO3AbFjp8627QAd4HtF+ke8cYtR+Yp7P7L9sN57qllbbEr3RoEshmdWI
kACq3tZqsthLW5UuAIFKVd8VBw2o9tRY570zHqBvkC9WtJllShCvvklS3jzk9PkdrGeFgTTQswzM
Cdye6V0oqbUa+R/suT6YcmE4/45iYWSh5UgB3v1CGCzbAWhXPghuk6yuOqsD77/ceE+uZ2nN/83+
CnuTKlx9qpxbmIc6Bf6p8qozi43hP4roqKSHd7wu7vpGl5Onw0N+kg46p0e3k8grNW4ZLwy1zucr
W5Izt+EUb76cRS3XUGQTE4gR3Jnfc3sAfca9+Gff1tL98fSrEZ/8TfMp6aPDScutvy/nyPI0Sz7h
QgdgiRS4YuEAx417NDU4SGVwYRIEa0xk429RuDvvmuy13kPuGTcrA32rKCeB2nzMryXp/o3dx28G
yQ29DICF92kZj9DqEcs/2bI8fJ3SreolMrofySfOhL4ckumh0GqvZmEGAyAH/YFvLxEq40+6CvOR
cvuhAxbnKRrXUcAM9XAOy3HF8NJzrXN/6OA88EH5gwyptOfRnnj0ygo5ISpzmPjHUwsmVBtvrhUo
DTRPPZ0Y8gqY0o7UOidC++A7m5OhIrVYm3KD3Vj8ow3Z/2Y5/wAMCpvfH3JwagMdyE46QEk/LqMj
PPIU+4EWheaP7x4Q069zxsmlTub5AD+YuLXyTd4ZOOkvZcNK8DiDcG4ekjKqKLC5vVtZy8Da9eKP
ATpbtr0Z8WxHWIU+aKVnNXL+D8hbw5y3pHy8gCNrvYQbhYYNX8qQLAokkufMdNvBOK6Or8Og6aDO
8I6NiD9vSsEqrIjee+eB9Tmr/Oyx2EDLupK9euLI/LG36OzlsbNrHfThQEvRVTqCGk5Np89DgARV
PNDtLaWctwf2ZZ59d3cVCl0KXpTN1MfamPGrvl09ItY/7TT4Iac09MmW5WaHwQu2fEqogg0lq/SR
BG01ldDR+Vo5dOltndWxvzeVrSJQRDiTa0qMBvcQ1deQvcIZJoHKHDz9XBbRlBQCMzlzVCfqvLE8
T+zy0MUENzlgJ0Q7LFDTZtYVTdPC3oQZceo8BvFVdPqgof34+trtrLsRCYVSNQ4gOw5amTe+ylaa
bKZ1NGabNQUMpp/lxULxvRl1ionJOXfAW/Fz3y0WwuPmcMkkgsTA9OzHCIOwe7zUj2VXJf+2clD3
Dn/ZacGtfhkbqJm0/eeeptKFlcfOVX4vJsI8TOtYizOyKqX+/nrRjzqpQOap+BRpoZ9dz2uPAv3g
nK0ue8Ne6Es3daIgJoywnoJO+OJb016+58/YfR9WhLn2eN87r1UOGY1C30tEgVZ0WPzYtB//f3SH
4iHT0lzQ02DT/YCgXVRIRLsDS109Wa0ek31rKQKot4/o7BO+Y44Nw1frfLxTgSpzZQx8+PJh80/W
J+otyQwJhJwA8BJdF/oW1FEnwMcNW52SVVubDwLFhU7S/hyFg5kVyzhJoiucYagbQkwtecTI9gQt
tTrfQl8HViAymfplEC0Dj4lbo+/17oFemLa3N8rfu2GsE5V+WyBVOsxnkq2c7n4iguvShOE3pKm8
FHv9+/bdEIqMA091aDKnZoeWKBPkJmp0PK5c9mKbjVP82CFJ9IfTq3ko88ZyfcGyXZIxt7Vttw/O
GmLYkwAJ64Ea/yojHtucJLe2QtHCe5rg51WACx7VVGkvJJTAyRNdK7ygRmvLVB+vWBuaAN8hQSs7
N400F+ERVCK0U9ApRdUYrT1nVJlT/HYdP0Z/mQbDKcwtJH0cPIRGvJxWSNoqEQOsZ+KmTBr+dcUq
WKqvU+xThq0rq+McPoChwdPOPkOi1wGzx/ZWpAX9jKAscBNMfngpFh106HcP4oPnqDRJKnuv54Cl
YwaLbfy9jwQonO8sItu49lb5LlSZxuZAdnqj5G5GoqbQivaArwL8CtRuhoczhDlNgk+sCXdGlg6c
KtXaPx37E5HOiKUsbT8v9BD6g5tk4Rlso0eNAX09UY6ZSqVJF1MZvce8EaqdNdqn+h8aVGvWtT0w
GS0wIHD+I4Y2Zo0YKHejjRMeMq+T5yg0mawmck+B9kHv3jGC6Ry/ihT9BcA4tuwOQx/oYrgVTguL
/pjIznqyATsao1YAqs6L3axVJWnHCroib0/JaFlxc0qjF0rU132CzWiv9ulkwoszSKvdBDKd0HuL
l5V37u2g2xP/8vGRyj73POr53GoB4Yq1/c7qZZCADP/f9YpKbLn69LfmrERU9pSY8HyOOtzEM1tN
CsGxeNMocq83uv8JiTPKolj4S/T6czNT+a9uISHhjK9zJDIAbjQ5qrQAvsMnWjwxn2a9xs0UItJy
XAD8z3lGZ2x3ug3ylPHnzrvUieskdt9fzA/CGQnxoX6sjdp2gnBSxUP10jYAquuTizeaaRVrhKNy
J60bQljqTpdP6h/yJVEx8zmZP1ECIQPFxHV6u73qiFQA8KeYBPV5gBo1Br6Ur+59nNTqOqEn5IQc
i7WAGUrlOOSo96bWn+KzqUGenL4MWxIrOI7PcIgpjTzl/plDUi6J3HBwZn2poU1nYiqAxer+1YxR
b4MxHCEoZCwQAnUuMWYdseJPDF2IzhtyS/Z5V2KJtNpQWs+dtvoY7/eDRCClnTN9O8a4TNR19JVs
/pmi09yPWfY+OV0dPe9bFRBNJYYhm+rLdYhHxwwvFLrn965YjMCIvYTyGTxYNsuAXc0mpeNv6ZaL
UvN4IDl8qGRwy+wNyd4EmiSRNhOaT1qWutx11yE+w0bMikYfLxsxz/Cw5LKBM3ThZNnr/cEignga
RhAqH7OHtNWuBp9szC/XZLW72lxSP65OQihixDDSGqhN7FcFQqbUZkMVHkjRUzLXhl0cvhAa/4LF
krOjHKue3lZtN59sTgswZtWJ0GuDE03W4JIldRtljYODW8jR4L4z/N+SDQM1P9hSlYwlLnRmEqu6
CiGK0mW9T0om6MU7EFXx67OtcVvzFxDVCZ1PS+6aftVHmj/dXVP4RuxXdAc3x0ViSpQLDIM/gG/W
b0fEBD+PgUOsj+5mIch1tYPQTuzMJL1pUmRzSmzAsJy48VEy8xcWaBNrCQPFosvheivu2SBbL19R
DAFrv4qfH/Fwlh9G/ltY8izL0ELehIISkvI18eL8wUior9PxbFjGCbI4YT0b7LEzTr4CCYvhKX25
N9ikr1fCCKEANoarzuFJxOFthay/M4n1A24SASJwOKEAnGj9EDekLSck2/ab9udizljsvsg7h9dv
zLCohhL/OuvLJGGkEigmrR8CUwds1wxp2s0iWrSK2yTobgieIe91wqsRqH0mjZ4gZxGajPywAN/c
/uRl+bk1U8ZJn0SVVQscIcbv/afh1r3py9BB8nkFriYT58mIuuJZOn3SHjhdgTBQDDVM4iD5owWZ
QYbJoXmu43ulrw7FXmX358GNkMB6G1PUVCEKSEJ0zqfg+2kuFwiq0X7WEuFo7dmLUH77MjilPjhO
74JvFGmvVYYiAiOLYYyh5c7fysfk4PKGGdqm/v5n/dJK+6atXhtNphgxKW6nJKuinz58EiYC09Fn
A4M2fdGkhXVwEp1ek2blfApkgfmtspl1TKvu84FO78h1d7awNFbXicfs3D3a/gIoqU6v04CvFUcc
FlNcqQ1QSFhgmdbl+2xpgvqNaYkFbyezXKe3Jgb8zIISd/O5QXLUz4j9q+CgjR15bOCAyDVV3wW+
XdsNn/KOIdeeOyexSaHaqMb5ZZNI5YuhfiZGm0yJ55nnLgHEbjqrg6ANvsKyGUG8cIQSiUEeav7T
J2lZcrM4Ldgv5Ln4sF3xrcBQjQoTF04MLtRvBoV8mUO4o3VtuVfWcAm93Z4ROV6sLelR5v7Kxol6
ChhTVv5O3TpMI+EtWwzTnQxYst9fXuM2niKmWa8I9sqZ4Vl0VZfyG8dgNidTyNb0oFK2FoDw/gR7
FrqdC9LYJ/Frh5Cx0L+SkpNF0jjzbCAjuy+sz5s3lHlnSeNwWu19lL1ZPAIYsNjxb+7r1wfzb2z0
W6Cc7pCIzrG1wwfyyRChHnJct7QDqQxLY50Xif2utmdBbKy+4cSNBl9drsrnE6TxjNo6vXCFJ63L
s6NnFsPfwhoBEzdvNqJqFFdvoyGQoZUTKoOWSUoXrlz3fiZJa00eM170P2AWUjdLb4XU96m7X3u6
3t/Vma8YQ0zVe/MOj48LGS+/UsO5WHfUUueBGXY3WuxYjMpa89RGwU5belyUWsF6KEQGWZtMEFoy
rMat8tmJtL1+43mCQhSUr2HKGRFfeGkqW/MlCVJ9ibX7l8GQbDIYKLTQSfJuGZdwLEU6SZTmpFkx
ljmOFoKr1ptJvHCW4AyEYM5bwPo9kkANgZ+hWFs1WjW2tq94fs2dEJSM5OIhURYqdO5VhXNJ4cCX
J94JqVn1MSYDDrMcXJl7kylWig5Oq03POskaVXgX8LwPAjp+wIlQJ2KT0t8ym6/Kf6//iYlsG2wz
fyZ68N5RQ62iTdDI65hIszPtPJk0le7r1Tx+6/LZFEtJ/mrCI1x0TimzTkbhy+3e5kAGVNe3eYve
6sqTJXzr4Kc4FIFqZz4FYSHMtg44nBLTKTJzuIUyQroX82vfwXDyjruPk9zEn9d2hlL5nZWzUHUF
tV89hpOsX1pddflIRPa9Qh4TfUTsGD7s8SJC5uj1x+O6MLmYwmvLDrwyEvGtMGMVZbjiqG0QwX2g
xJc8Id/yV+UJbAzieykcO630PY3b9qvQTMAX8qrYplYw/Hy0d2dHodxxE6mxoaHV6zSVUxt3wJ8U
6AqlB2zA3ph7xcU3Wfh1pLMLP6+5RKYbCkUs8gL37QbmxFw2OjApie3N1Bqlln4OLl1y0XMvzmVP
wO9f6yPhbwsrSHdoHjRQWmY/FM0KRyV+SkFqs5lBRvB049JJpnVnkQpfOfrzXxldmtxx8QHUzSSx
5bn6XcERch3y02aoxOkCVQVgN/xj4B/Tj8ivS8lUlCnv0rPCNfICoYTSYz0c+c6q3uFrTvwsw7KM
Gv2MsHZvxbLzjmnUTKioFbaSZPxdYYLgXKPGY4/VcLzNSqTsJn0LW8hghzQnLgqxBb9IORUSpG4e
iGn2YUM26CZAoY1QNrxwqUI9ckRxcjA+gpMcK9ERBvnq1KEzXATL9fRxI986rNJMSoJb42HfGywp
TmOXd8NP31rZk5obRiHFuHFCDs2qmhDxCW2u/GAbLc1RLB+FvKkn6U2yK5TnBBEIZlLafR2Jr9VQ
xSuPs+nXD3ZZOVSmhNa/nA2OFkpCap2ZPpYOqYSxBEs5NDf2YX63lQrs/Trd9cP4nFV0ed6iJ+dS
0CxTeJYyHUEk7eqg77ePBoRjTHPuxQKvrUoWdKH3Ur8BrxNzLp3eUQTBbar2IXa101XVTyopqyaH
s+E+K5F+EmTB9IET8s6QnR8BP+2EMmK6ihw7uG7YAiogCwPD7Zs9lxCW8vmSe/NnVIzKcMEqtyfs
L3AfCSK84lRXAftUYv1yPdkMC99bAJRKWZ0mFAHZfT8+w0R/fKZtNIF4prgfc8sx5u/nfBI/GK+5
K1QDXr9waJ1BpI2XEzIpQDRIxTrD4w6r7vsD1eEMz7aZdoV1VIGmTXZ1eF3/rXapJLBGTdNfhR71
7gGp8dZOzf0k7TnbF9HOjzVOUUYcYKccDev1rAc5tYDiDtwex9A1kghoRBWNd75XZUuHQ3ghi8en
t5bXLpjUKIMLuCJFXVg/gC9kajgV5VLOpqyQeSXWomzrN2UL9kmP+66ypZ0rkEoo01ypbzblXzlS
XaCcOwysEiT9pYy+n9Nnh6Y/1+z/PxJCqEWKaY2IkxpYIWjE1o+e0ggw4eWvlHx1teeB/wke8vD0
UHDeGxwbpbzSua7u0/axwiVrbRGAhzM8ndntO9uMxjdQXrhDcF1uwMie0nXqYRVCJTvB5aVLUFpQ
RTIGOghshxlc0hsLnU07NcZvfb2DSdQ7ABZ1ujwqE4MmKIqcPfsgsP48XXKTsqVtxpxanJj/68Td
OPL7jlZBSpdELDvmJxPxLwAALb249P7QFCYk6Zra2mweu26iHvJnp5whUJZPyjUONqll6ie/Zb4+
fthYDl6oB/kak2KI01dNboZOw08b/Q7yPPeQbAqaHB8ov0YrCXmXSi6IopR5Z41O3Kx42k0Z9f2y
ovSPTAhRchC8YQFRDbXUjsXWoAsj6IJY2sebkEtp6GobD9eCTF8/K/LQ7nZvRVvdn0ptAX5G5Oo0
10CUzw1WDnrFSThStGcxMDAtRqqSBHuxbCCp6Cwh0R133lMHkWnsqdyMATDwmzpfOeUmE6uF7mBv
iQNJn7qUdXee2ZbfiSohTqYloaXOO9ByzND5R0wMPTMWqSqRr/02t4Dx1YYzAuEN+uFeZOg/ac4C
7++FcjMIIUgtC2QRgnACYMwdvQsi2awZ3sPrLjQL7RpTwhVvqBSWDX/8fK5xWTfSyhno7NBUukv1
T1TlASE7vuAFalosHmHvb8v5ALQSO4P8XP4aT05pW1Fjed39qK8fEyx33B5S07IuXkTsJ+wHSoWt
LfltP1CqqQniw3WHTG+Qcw7yH2JUr8Me91sD3vYQ6GbzTzRKW8zwQtLuRinzOErONmVI4x0v3YMl
QH23EgGiL4E3PH4P3PdSMyXAjsyu7eeaT8kzvAcUdG/JxVRkXUnLWhKkGsC/Ag7pmXGxeOYzumS2
li5NeDaFQsN5lvAKb84t4Zi7Cj/qyN0NoTEeqKlGZ9jij3WbxUGp5wv0H8HFxdZcXtQdX3GqzgyP
hwhZGES4l/kRTjOaNHDJ4Kgh2fldfXoGOR/cRYynW4ci63/hinew0c7tjVYjX3lupbe2SlxGdrT0
WHS5nhgQT1QgmABubm6LAkZRgdQEuW9Ixzqo8ss+FpKWyHNtfO1jMzdf56EmF/itYq7/k3l1z7C8
6F1QF7+z2TKyG1Z6N6aaxYULRskFdcbmzb6mefv6eoK25aolXM/85JefcrIJqrn6zrMHpJTUDjek
XvkdEEmxXmppMCxMwEJISo9CTBz4S+CuhCQHFX6ynyJowpd7aFj2n6FGqedMW137Uf+pjR/DoQqd
VRtwF7gMgIMdJWI7Uimw3hc6Q9s+BAVd5S0KQC1a+zpmJM2MRnMuhS6wzMZ95YpU1yMuxlFoP5at
sdxv4FyK00wtFA+1ZbGPsKEaO9GctJs4+koHNLT/dOpauoy0elunZDiSoVvm6oTZcW4w9mQCdhgY
7/xE0SNnow8dxdC+5yDjmWhRYxUckkXKNS2zD64hU4prG3YJprfS6/O+OaXsVJFM3P4KN6Dm/hLi
KG7uKzZ/r87+VVQNYhXn5GBoMAkmx9iE6b8uUGoroGsIW32B9vi4cBYks956EnnST0j5TzYBff8p
KwkB1jksz0OcPW1Uj8ZlIzsc7D5t2GUdrZi8zimjq3Qtgg/4Kf5OR+jP39C85gB3WWkZlR8XO799
hi5ASlhzet95lUPwVKOac8dEINWyxDWMG+z0RV72Em2G9FEDg3zAZJJFQ0bIZN3ZLVojOLQJYHAF
xKMxKJU015h4U1ZRFDVfS2iIKE6Lg7tVJOSVASMFC7IT6dYtfQueS8I3N4ZxnaQJFcSTiio3sOWv
PSStlelC1ujo962PU+VO+2D9nUi2NCNcSk5171mfxOTmwa0fTVLLlUqFYnvXweonbZEad5IZZl7w
bRoHdtcp+1bJXzitvgD5SRWdhRDh7Iiu2icQdIIT3WoWgwgFtBxx0KH+l8nSOV/xpEzgmRWD6PR1
1gDMGcyK7jsn1OPPjbgPTPpHfkx+MNJ/5yUT/SYcAsL2w00hD6hgi8xGhpzLlgSkuZZqrK+uagiM
nUIYgqH329gaFG+GTYg1EWcQ78yzV/Lf3tyvbmakybhzKQ3fgC0Ju+7yHq46sQ7eDV9jp93JU2ZV
Kf8W7KsTtjl9Zo2n6zELkqPUlT/MLDi9qRfRDRjAnE3JdaLh37ofIP/Pu8EBjcqzhPP7sgXnOfG4
cN5sW6fIDP++EM3oLghCDovKHxCt6xZ+wanZILWpESSg81ANKCy6HVpzT50g1xvaFT8IFje5SgZ+
La2D+jauGAHPEFani2tifS8K/6tTa9EZmMNoGonv8xDLlyyGmk0Yurkjrz6K6kOTRPGFPri4Z4J5
G1HSxmDewBoJ+mMEvVBaECh1cZJ87EwyYtAAuYDFLW+Nou7PAOJApOu9nkBP1ddv5VJomUL+iCYF
EZn7sTLn1wb4rzf7kiieKrSi8dAxIgw968U6RFUAoRnjhxb26qUln+eGB3/2Mkr+aFLc63xrZHeQ
JJgZoI3tGqoQsOWT44+oHLZSpnWgGnS49cy78Vjk8SP/d5pKVMdVlrVZxEd8wDlqIIOIdiR/Y5hA
MhL0G982GEo3uDRxylkBlOCFtW3ldk/FSaNzQJXxMgxGlRh2K2tMZkYAplyAL8rNyz6kCJT7B8Cz
3TScjrfY1xlLDxkajnbcvR66JSOsH1Za44Y4AlaLRSie9j5aapx7ypAqUmtK1OjwQnvhpw0fcs17
6lpd6vKX69APZXwoPFwvHPqP9U1+KRVv/j+UzjS1xq1e0hUMnBbmj0HPgP+X96VJhlE8e1beIYrp
lNh092vTSNlBg0ncEMqASdFWqHBbnd08jJYKNR2nxK5kExgnSYCZZ+xAQZDZmQa8EaN04Rlz9EJg
v4hFKjiB4A/JHc5xongaKZrHFsO4hDXNywxPPOc6G3nCiAYnY/2hKFtPs0STWvVo+H1Z/t/jAX4W
xdGVZdEBPZBPMXbtbKsG5EJmk13uGSShkN8es8bpRTwCts9hMpxZ2nDgA0pPRR7ap+xBo8IZPZ4y
SHmu1SedLAFPGB7+qgLfUXz/n8/CDC4rW2Mh+mQNw503UElHuXnHanisMFJSCUZTT+rCN8Uhf641
hUu2IBhA40X6teQGMLc1k3nD+90gJeBY2o8XUQxjePA3yokebVSEjRBA0T0qRHvERMLMChbXJL4D
IuKOJQCKt0GTbYqfvZBe9zbUHxND7GUF3O9ynQYzStaeFqCHeshcx7A6O95e1yqyjuHb7jVjM2Rg
OvHbnFiFq0ZzyE/xMBC0s7B0YAkxEew9dhtl7xF0u2ccFtvXMFpdhj9IyVpMIDlPBfsc83sMk7aw
PAe8885/8NrofiMqHB7E5Ww3Qzo/qxcoSZOp0mfWm0uBcLzOETCvk60SPkSWkxqKw97lDK8s2Rpn
pZmwWY7f6vdpT++BLglN5T6cU94t96UQOv6kXDlc5QHS5ZQ2TquopgISIuup6JuUyiyx9o+KLLeD
RGDwqYa2M3rPpf9wFjzC1iGHJdl6ukNVQLIoFM44HNwWQBEEVea5zzkZfX+df3eev0zKFNqyWHui
11zSCgvmxBryEdxz2tUjDVCYQ5PqM+eY6s/eOfrtq3EGEL5TD+dsXNrKyP68UePWmfY5Hp4ZhVcY
QLAfywuDmqtlzehRCqhi38TNpRG6berwgNZcrNfEp7Ut0r+QlwY+6HBWK5HAyKK/jr/f9D3lKTxQ
pO/vAdDz97Ux3gfU4+OMagcwbGqqcDajhhbWa4usB1O0Gczw3DAvCwFqS2ApwEdtCKUjFoB9OK0f
wYm92U6dedgtEVZyfvWrOF415grMQAfLzgTeKSjVPCN9tDB67ka2tk9IHclSHZJ0rBf/Izpeorg4
ox1ac/McWMAiDn1QbcEzi6cb5sA6Ax9+ruibJDA+t3jqaE0zgTLy8LdrG1vFhR8y31ar5DBETUYW
kZnGNeK5npTZ7h3/VtGUVdRlwADPVRelXciXDEixMO5I+h2VE88pxYJ7OUfHYGJL8W4sm9zVqSCS
8xOf5AuhsCG/2Yu6QQYAgNNS+4cpvx/LHjwMlfwqbnvwETKhDRWHkvMi3utYpVSQgHC/75hQRpgO
mBfGm/aAkw1vQEPJvRjQ6msnMwl9qiMMr6o1F5RXv93DUH1gvuve5u/NFE/ppE+Uug3W8jhsN5rA
Hkewy8vFY/RqjLdwPVFwScguaHjmUMTBO/kk5DRDDWKuaH+JdoCN4tlFnr24Y8bTtpoW+Z0y9tDw
npuHRxCOkd6Q1IxFtaGQE1enByV/nMmG4jVYugKvDFBW5d7/PByRIVNkf7ZfcPdJ3YR06Rznf0l1
re7ogEwjdriHfkPuxoBmXmZm/7wG91NJBLwu/+mEpK62YkQucmnkO7/HPjYGc1FgOF6bliPfmDaj
Er8WIRn3yncFpQOQxySP5LLL6Zcp5AqwY2u2XNbjlvf665lrRdrXipzeNJNpW/dxNAy+abrZW192
Y2H8yqoWx1pbGY6t3MFKbHA92eNhFm2HpL12eCbWPxlQvVKAqAgatkk4pCKB5pYmOLaZWRtDVERX
S6Wj8j9lMXUEt329jzVGqHfdjBdi39J+jrLSGQCuLuP0Z6CUU12mdOCnjbOu7Js8sM8EjnbY+jsz
eFUqATkkImmipgQyFYdtvhy4+CWJpuowrxLlvKQls9EqeyPNyLAJPsvIw3Y+RNXs67QShONxCIc2
XrQij9TXN0mzpvVKQZO7atiMU07oR6Ral7A48QVDaKE5iAcFvOdzG9JjcQZhus84keXauBowN2wy
QFa4obwj/QyqkfT8TSWanGDl3b766L+cvpczMRh/Yhn84i08w+kiHYLrrzud8tATqE4a4NuvS4yH
kq0QaudLk5J0YQuT81jDRea6oNX5MyqGk9m//3x/Eqk7NgB5dGDVf6AUMhPomwuYqQWSBZumdsLT
DVTM7v8ZJFlHznfWKLl/IoYF1YkqS/XKiHRhzLgKhAKsWcFXCmDL6JH55fLz7rhjKZMZVmmgXwfl
CbbHuYr0qSFc6gAbeG62133kkBfAywEP5TzCKAcwl4w1jyzM0MOemZXPTyocI+qG0RH4Du1W6+cN
7cc7gHjDpN8h2F9DhdC8+wCGjNAaIT0cRZFx1Hh7CyvTFzAaH7SnTz+bMViu7PZqVAPgJbGzU9nE
ydfSejEODd8dFTX5OvdtWlLfx029K7+mzQUWzvTUKd/vO8h6qq1kooifX/baoGtPnX5qycnBEtvL
RPyQOy29tAipoU7u/V+v21qY3Hw4hYUk7bRr4wKRM+bFvqkwnYdlKIUmngBnxjzzMpBE12C/Mwh9
aQphWHObLz7bKKe4t5wqIMqXEyOsi/l5YgQiCZL5OOTlq5ftecDfpm20g/BW4ZX33lOzEkXhFaYz
UuPETQBLt/vFWAJGnwft0XwoELg/uTDuEXEoTrdha55IQZkQh2PnYEeOxVfWnUl6LRlDAbB9DoDS
y8y/qXp/oCVYNyd1Z4+MSJY/0cGTU3SsAIJ24mAYw08CzlYe5ztcI5SV4g6g2Y6GG2asOky8qZ7l
iV0rJoCepWSysoKC3Jow0X6UD+PRyi7QpEekcc+ERwjS5tWhhc7tUAKNrht+VUUdo3HAcS2ZNeLI
ZaZuk6yYEYhMm7jSFnNN5eITuEvZw9nZW5DrtLbjGLYxjZujos9jJ3hkjAE3Hmf4qa63zlcKYGqJ
MJUD68hQRb1Dxwl2lmohmIc1EZ4uFOrBc6QbO9rq5P90BT2FRj/ATCgLiOjuycpEahXkCGvofZcI
JkmLF7OL4bjfNQuMddwpmLG3Pg68sG3Wnh7g57W6Lsdbm/Ave7nk577O6mweVHCMP8jQ3/q81qM1
0I8+eFsQZC1om8pGf3uIw64hqzv87VodAl+8RHQEo8nde+GALLxlPPksG0H2EHUFTXLIIwrzZ8Dn
4tBQ/deErcseA0CtN5a+KOVofexsZaYArYmG9nkfpVsQrtNK3/rKJClT/Kf1AZ+Zuw902aRKY9wM
oJFM1bFOKi04hJJ40232n+gpkcKCF5eFgQvnYPVJNyD2765CeX8kZ5flY9b6OpFTZm15u96IQ9Ty
tD6vZ4zb8RxYC7MsMrUAfP9jbiAmbKCDvspEn7RGZ181LQY1LH7/OCSa0kYG6HZ6StUkrMHuWDzS
iUpjPd6+NcYbIDl8H/pvV6dD4QtafmN6WtH3WhHgGRl1I9rquCXq7CaKPzi1K/c6fsuO8KNNFwnt
MAsc2+fbRqz4BwzjXNTmVH//HkMfladiHNiczs/dppP4ZxXzM7LqqbcyNOcoS1c6C1JS4RParIU+
ZpaNpkCRqBUpZuvKR/ZlDALiyAyOBBnOh4NoLuW7sgtvpa61xTWkMBQ8sqb9toa77EsYdayIbzDH
Dyzd9ntVZVoq4Ay/4U6hQaRRofRCP7/An5HxSiShkxnXv5zhxuPnwVG5SdKOta3DDhYDSN0y9Zbf
t3bxgdEhBXR6QoTA06dHooLvyCdabwxIyEv5IPISriHgWzYKEBelmR7v+vU51IXgpFe+YwBMNVW2
feDyIMwlZDNFqbADpxLv6s0JUFchGEbhHPEy3v5FpgLu9IxIG2++2OaQ3IBMPTuXlVgIv3V2HirF
M7fOlW3cSHMMIkY6hzRWxct4CnHCMjhGroDwDPgfTMLUg5zhIVEklkADuDUJYtdN0S+UXwvPnTtD
5pg+tpSo/ydqX9JxWjIgND4O48wJ2UnDahuob/kkmFDoLUsSsUEE5nSdcE1V/ShorF2qjSlOKkGy
xJUeLXzxeKrRitoC0rgzbDFRWSQd1BerQTQ8nSAtU97NJYBmEGk0Xkd0KnscJBXJ6lnojfNcDLKl
a7jM3NaSa6WZOVkHjiKYnBigIJ2IYGl55WjMLQW4zGrVxAC0yMHhyuzNZIlslXK0gAeWp8jbMxor
skXZUNZngVVvoPP8vbs57EWjI5DTSKlufq9hUTE+JmKZqobPRxju+6ThyBHZW0NcUHdQY+iJ9mtg
dpFDiLDQ7Ltq6BVQCAh31X0/cK6sgVNHcsIPub6VVaBGQHORe8WpQDpBQdTSAtPVdbGC+Hae5nN3
ddilA0vfoEE2vzmEDt8jy9Hj6zW4LjH7qhyqsLQnYhG1f9Bbh0LvAf2JfCztuxN4EiJi23/Nn/0d
bedlIAFOey6rjdx6QXFlLFfxwn2F4jhglRjfHpO5aMaQkrsxqzYmNe70OgFzbcBZduwTHqOjokHz
uKt3psN1pCBpw37HMLLhKGb1tLdG3Pm26LawzQQz8/HEeca38Hs2aQHskxvB00KQ9bPUcXVoHjv8
jW3NhuIAnvcuiB4Gr4MP0JiSLO8BOmim4+PIo+iDN7ese6hCU7cxAg0vaCzD2vuHsFbTr1CqLDGF
nrdVYxKm3K9f2qTbF6l8Qcp462p8rt0qtmp5PKvOloF+EX+vgXMHaTPV/5aHfr9omWju5gKhI4Uu
6ICQKJT0jTEmgSmA6+1wnm+o1nX/OzaiF3BFlTqsZP/LcJQsUJSJT9Y6mEUVQdqjoqW4i5e1henG
flKTn3+uPGzEmDQyf4E9i72Q/wRyjsBQG7JTMVWInNw8/QScPRMcGYDQH3RD8N139snSfTOn+omJ
wZDpZrQG3Sj5GPz7QMJvaL0M5fLq+Ody/8QM6r+FCipm+mzRv5ONF4GrdoqwaRnnL67fGs+OzpUC
E4dXRJwhA0I0GKhoPh4Y5b7wVE+tr8ErBgqZJ3JVSENJN9IUnrBwTF/99imOV1i8Tmgk42xK3GQ+
Tv9jm1eVcXZnOLKrut/KtTdqvsIw5S47uPHxlt5f0MzGSrfVCKGfTmTJ1S6tI/0DylG+V5UsGK8O
ZeOe/Vup4y83XYeyPlSRoEwnUrHFL4Z9Flu41WS2GMeo+YqyXHWlvGJzaK+kpLBW1QUx8wn7VgGB
C1sbz/f3WP4z/NYuwUeF59KOP/twhCrIQr+GXSqV/o+pBBhh3cHwZL3yHKLFMM/cBG6QsVr3rL36
+0UNQJdrWUE51XHcf4OJKbqmiDGFm3qWCics2Ik5PcKOf4DrMHTZqX3Pzjm86wVOLLzrfkQcEkfS
RcSUhnQCF5hzL3bRE6Lo6jhtfyVJ/1SzHRQTqFbWBgRmEE6mV4movK2pWEhbodLtWd0hx5esDkzq
arV+uJfWdosLA1CnDamfTC3HK5OjfUtLsH89THAkbJje88uWYmOe3lztFnXgQbvXa4UKddpf0pz5
AbWKYNEcEJ5kZn5GY8do0rw0oRO2ylj6k6Hd4Hhzkvg1bgBEm5vkWjL0H8HM1zV5CwGBfTcgEBxC
n3/+pssSifPDnaiKaJQD/hk/8NzWT8GlosXbDtmr2APUkYMiUDcRlgPMtPRlHbMkdLZqsftaA7Qi
iu4tAwJ2jIlZzBgZDwaMn6fPxkOKVzJoVmn+lpJVWhnh64hlPJxWLAAaQ7QSPecvoQ/sbo3N5i16
hCnbHUv6ObZss/Sd/R9EpPjdOLd0aGtufitMloedE/DVSg5Fwp1cXhsYhpF3vwyT3nzb4di/p9S3
qAGQSY3UIpn2DlMOvrxJVJZuR/GAvRGYO6YIy8A0jVyIOatHsElqBXZeI1H551Q0qCW369lM1uIb
XskQY30BDH8u3PHXwY1ujGR5krL4yr735qq/q7y13Yk9JGaDcGto3bmxXHDYkCXTtwbXIA4tlo+a
RdUfSwf8A4AqG4ryFS4Lj37B2mlaOd0FyyEsIur5oFPmnYjSnAvbdmW8MgmCkt2ufta8aOIwT5IY
GAlrjDkLNg8o20yUck5ND0grIjS6pdKyNaIFoKdEOGYPh4nSyY9nqQ20vsTmbGG4VSDY36xMoP8H
V5SabtdZaZjIrUdkSsuzCKL7H8+8y4Kefh+e0HUjzExziwO8xqQ0msHz5xLujSwpeyXpYr5A6go9
ilPeXQuK+SkALBqxy4srOTrh1/Kw/HVkHKIEkfkRpgU/4f6mnsvaK1AMAj9S9Jjt3LJmypu03+sr
DqUwz/odH53VC0ynB5oGBLrMGfp3flRznBV7qRuqP/aTtkxJ+tLb/5ulMBhDv9Qp8IbZ1CkPAcDn
xRzR5JwxcDWC4wNhrryw/EYyQ5qRSpQ32Gt9T6BfhVxXcc9ZwnFzUCrlDX8hZwAiHqmj0FAfk2P7
n7RpRSn4dwFoxdIqCXu2NmsezXvlgPM+eymzNzpJRazXmxhiJXLLQ/lGzu5zsWn1ENlw93gQY9ZN
IcEPhYSOa40Fyh/yoTpD8TGi34U/mB574n8GMmOSsI99urRWaTfiKif5TdbY/WQ41FhqhPs10DSO
ym0W125PviZls7uadrbAL6sTbCWj3V/qihmP8ABdT9adzpuDL/BOhapzsNLUszkxo3PcXYNUl6f+
gSz+xx70CoaGpjN7c32CLQILowRVdko6mJJLwzvynHfmztz2vxEOBitR8/9s6NwtV36T9+AgawQr
2VMdxN2Xdl8cd+HtoTdfIzjDoV3S+dTow9Gkx25hTlGn8hu3sBPy4CXBjNSa9nL2wdnWH8LUesC1
yqoqSAt9H6oCrQLMcIDqeXaYBbyQZ+mV+pecKkpZhlNX2WO5tFxpX8WFYEucsF6JxzJLPqpcRZqy
/CaeARmy3sYzvEOLambe0mINw7BUlLizdi+IDty73XV55zkYOYsgApo2kVJku1Yd5+vo80rcNIoq
PJS2N3lHKBpkQpVKiBSMOjHLcpE9tnZqZcje5H6xCvgSg1Dl+O18FCklCopyWhTHFh62n0XeK+Sz
bESYJddL/OrjPbckqTVjSu31uJH79ixuzd8qzxhefLsYCcXj92mMjCQtIN8tesEt6fbCH7aFl1lJ
cEbR56HoV1d/GZYGY41rRj6SQ9Jdb4mIYmTcP5SSlMSpzjQafMTR0DVjneQnctLSCJUcyHzJ6Mhi
W7rDmD3yeQ62No4kSUNFn6E125Dqjjzw5ciLC4p922OJSdTdXy0IEIdB2CCmRDUryI8x5xie7gVo
buwA5c09grI6x4/qitNBj4lCxmKa/dJ2uQLDIn4ymSirgCVQ68EEs5olX2dfH3QjJA5AfYm4SoTF
UAQDm+/u9jDok28neKhsTW1eGmQqReqRb/hPKsosgRCp3yGtXteFxuLLO+i40CH2+sWJzarzPPpS
f4Fa9oxlYqTQcJ7xhPoDdEqq5SXWF4I++nqAZuF8t9+R+VvcE9wIkObBMqHueY9VYQJbzdHby5Oz
QZ8Ct4mlwalMnaQ8nsul9/j+2ORTQWAa7pRjRWl1C9rQ14HMLSrjZi3DAA3oC1wiNBOK2XGsSP0q
3x4c0PVmvFJ+tPHonsSOqJt9tRT+tPISWYDZA8elLfAaOuB2joTOz2KeZxfEhFaObUB6OHf3ZmLS
8Jtou29UMMn2nauzfPDyWjRRqiDgv4J0COI4XPp9G9CIJzVLVrlT7BIOXQoAbc41CUoTweIik97q
qGBF9LEZiy55Bko5IPM5je0bnXNxqqGaR7tecxpaPOVZ+iQyBHg40Ef++wPm3PiPE2uQbs9P7Oox
dUN/JMIMZS1hktrmomazKRhTKEAaRaWvA3rCvkqd8ZxG/HG7wTZ0ARYtD5okn2KHz60g9SJ4qIcu
oyBLVA9/1D53r1DnCCkKkaia0vXiiAbK3pBHVZ7p2xsYo1RCNAzYW4K970k5PqaBiMl4Bs3IWjMj
15rBZ9HKZ3EdnbaYZmWHB9GActlzeUpdfdgbf3nCmLnGVlNh3kNJvBhs4imT/wh8juNtY6KDeBKq
YRZGz/GH+YQpNv2YDrNNNwa3GbPARkrsT8zL0y7MyyeFAP0eKlYL+0VQn9bWe6IkOVQ+hA6JtqBk
YY7QMabzFF7papTkkWoXObH5Vj4KC/Bb4xVgfPTcuPLFXGpedgaDZMKBlsJEzvVWs7CzwBbD8fLU
480LKJJyQUUX5RgNYs6KdAumlDRf0epA1g9ePtiIn6bQCgVInL1RPv4kW3iF2HG5zbCGl8GWIVq3
pAsIi1gEQI9I17tMtM16YPlFso61voemXBtj1M5ErDUbsgbBIQHIcmQeDG1zFvzywzwJDLC1zMNw
GFDPB6alZfnoVSSqCz1C0XX5s+T6jxq19MXgCI+8i9/IHH0ocC0ntUkvfftvo1v9SJelAscUdDNu
12PA6BJ8GYzOGiHG5/ocOYPocLIiqusGRk3q4N2boaKt1k0tYNDaGgzskcOoBCAfxWXtjLKjzfw8
5yqPB/Qq1SuI3nmPEoqCJeWCcrQot3O7ppT0gpxWm5iwK3YbVE8w64gH2QvHUS11uJ4cFnk79j5d
mNu/4rF7qlW6dQJLGv0yHb2wig2UjEt5h+lGCoF0n1vVNdfaNg60rQjQVE/Td/16rrwN7hOPsWdD
crd5wSbG+zRTqFNv8mqLemgW6Uh3sci04Qz6kMiSruRnHBzDG2aaQsWsm6n2IEUwsYIdzV7rDHeu
akEkvpULnpi/VA4P/75omqX1FWzMq8xmCnIXfZjfsOZmEaGnNAMx1flJ3Pa2wZyew6kvxkEGZgyq
XsUf19/QKaM+RPESpBjqb96DVHXpP1ZwyxMZoHoNzLtRoOMBCGXNtROHHEoYBX7/J5ZfjTwhpSkE
zIqmzioPv1mFHe6KJc3rV5+tg9MLNfEVwM70ow8RH88QGaBqH21PgwDuKcYXkjeuo3mQPreekTou
vedT5gE7/gj55GWDzjsDSW9uagQIpFaEs1idrixysAWaWTvpDfWx9ALACWYIexaxZOu8z5fRpcVg
JNGkU6eeOIFlXsiNmURAOeiF+QQmy3DBwN01VpmEv3hP8JZromOW8VmtYt1BGAyeGg/sspKYxkWr
wLxAoWLGCmWIds4q88hQe1jsFvXicC6fP9RqVyNCsDALeGEFVAFlf/BPK/kj6iTAx+QkIloP7Gdq
lqZLqR1ZKGpdfxLfwt2XB+Zvx3Ee1GomrGf9wJKOVsnsV/W9bqUkhUtHF4yEK9aMIKR+fLxtWw12
I4LRWlKFCuvGv+Rm59jM8VNkLqnhCb7nV53ZZAfimTZeUO1aAven6fer1ENtpGe7gqyQy4AbJjd1
uP2Lavx20JVDArIsH9vcMhgGdzUzfVrinECxifR2jOs/CQu3dgaPGu0xY5pKn3Uj65KQxl4xZQRz
cM8aWZDw47HFbUWBTeX3sh7/eV4cvk8N4EzR0bYoLti8Tio9H2GX4Fq1mRfcvFbauUOj0Vo1KjNa
OYU1mxyFF3vKMXaMeNR/mAEC8aI2klZRXf6LMzjzrfJ6HVscSvZC65WO8WXv53WeI/K9pWGsYwNz
mBc2oeqXF/6c/Nvojh2S5z0qkRhh259M2vqB116XA1+QX4Yeg/ie4QxwxdyiQL6SoGdl3Vteqb1u
1zEQO6hDmafRAfOyI6MVLowT8yEcUucZFX59CnTtanWpBPm68naqcZreRizeADYO6pP3cpUzrkqx
e/I1yEUkysXU9zXbGJ6b8AsERr9UQnQygmyZZ01NZ5+S364vTzfYkwFyp5UxFYcvUOmi6C/khaK9
2Rn/i6Rqso1/OZ6XcJ1uX7Oirv3/bYc4V8uBxwn/NeJyLoMVyPcVfrtyLoIXvWPajRI7D5HG9a4T
rl9jt7ezqWOCPyLMkd2aKCS41aUAx82zm7fTO1bW1fPUCckaE2qvQUZFsoNrPVC32zbmKoDtkhGE
gRy+bABNMjssPxFl7dp26FpaBa07ZqEdC0YON6sZleFL81nS4CivV7tKxTWbnJgOA/73w7GGsK0s
L/34XcsF4U9mlnZsRHVYBIYhzXVT1K0LR65K0HRddKxqCxhVHBc4k+zPNPbn1HoiI1STi3/acEi8
ThEB0lyqzIK8K5Mm6ge+uw6atN60nhjtNUSaJP/aY7sgf/LItk4kAbEvNnAaw/hko49VZ9RSfUcB
pEBtHF+VK0IaC5N82BG9+uSsFgVOQw6E1l955x+suB+doKXae0GgfyWPPjntHWpUdlY7eivoouBh
V1fWkv+9AtiR0+3GndLphr4kE45dnBTMHFKVbkuWKNenDVjT+kqnigLPwuKmVBiThG4XroeJDJi9
YFn50ar9gNQWazpQt/+/90lbGzYo9AfkhOwKGsje97ArX7BU5ViEfOHydjVdaNkWQ/T6jgfOmkiK
hgo4928s6tn2Pxk+wpeRs/Vbod+T2jTRVMxyJkcsCcv+8ShCf81shrlb/93NOYv2WTAJZrUBZYFw
OdXakPmUEqJ2VPFFuH2eqBRfH/EtlS951yzAP34R54GcagEROsNuAqGfIlQvbk822wjN0lMbhkIr
yW4g2eZTBKDrJygwZfl0AxoBDjkQoGVWLsSGpUG/vcrGdi7QLWiuYOZ/Pj4I/womaqIMyZrOCgh/
1AYWCu3meVNCx7JuY5Y+oPRdtBSzI+glSbE78Ebjf5GxEclyR5FAuld66nfu2bCqEtL2UuVafDIf
WtcrbOT+OYqYEFF4L4Q+zm5Ticrrdwca1cPec1Vq+ULJn/OYZeLLauj9oI+BhpPGO9vY31rGVviz
P3whhHaJ5Ten6N6tY27IuBd4DzBmCzexWrLJ5Q+/8Ec9k0J8n2cjZ3ZBFeSnJPBpbho7MPpUbUXN
438dkl5I5cmSVgXLCGkue47G7T2PJvReW3f4QSJYLXtnsefG8GWVrekLQ5B3rNp/ynb48LUVnP7k
sM0uF/Hi8h6JCom5QTDCq0pbjgdgWCCbvLA9/Ji4wsUs44aar60pn98wkei7+rt9MTqUl5zQXSNz
HnGPUxYOz1l+c/JSHB6HXcscIVzwqnlSrt8Y588VED8/MxjKHq6fo1p/MYXI9/cNvduGHQcmzpWL
pZ83+VdsrafdvDHI1+SwlTcaMhtztSVtwjzBFbg57a3x7bM4HbdHlC8JMOKQFFjo6+pblzScc6s1
Ppj35CmNQ+SKARJ/+e0kAn/a7jjSLVBt/hwEPlRnyMK4T1Rg86KRsJwJuVTRWef2zxCP0HEW3HnD
0C36nhZBMlAdk8A0WiDgK865xC4honZnUeMxCLVj/dcK0Ear8lDVlFRrI0LW3poQR4blUdH2RH2b
+Ad416zfyKL51eTGMk3Z0F2M0TODdSt9TO8xuK81cHnwHBMbeQwnU2jzVa5st1IcMRPndWAjbtMS
fNQ28NorEIaRkHbJ7htq8qwPhpwBDoaTdEThLssY3mYdGmtEORLNY818TOeraOYbmcb9yBFmNSkR
WK1ro79GVME/QdYn4Fsb5LzzvKzt6hHGEeZjheq7h55/7cFKem0Ts5fJUpEGjV7KhesRpmI+5HMI
2JL7+yUEf1SswBc01WnTKJHW2nr7bPujpcxK+l9Q6++4bQe6R/MfEAJ3BxB8icQplaGvDOp56MxG
8xYeRbaDfvKE9CGudoPMVqzlGlzlAxDcc7Jl4MRB5dG7LHrR8G5RgUkZLrKBzvR8x+nna1Lwnpzm
wYqAqEhvo8xLOXXExqZ/2I4AT+xeI9yvYwLWyRQ0RRUeRAU0GCpQgrfU8RXJaaibkVk7FgKfZ70+
BJhxt9huSGs8T9If3Cs/BdyNM88Mu3jDuFI386+sDFZ6S7DWxQGkprcJ0x63lFrOI+9YFO3WHy2x
+sSsmV+QXBx9t6D1u2nXnndQHvRd1ncqV4/Boq07hC/6qXzqfduZen+Y0eWPZedI/8ZFBS0hrFYl
XXCoetvgRmdVtxd0VcjGH8Bra+P1uyP7Axa2J+Ve5OhSsiXAfXJbPyATEinnumwjgrHQ3HLN2/wc
ElEPrI9PVq8dR+kjKzmXaZMd7FdDDkucDCi+08RboZ3IdTOAYJPhuWlsIGdTi+tw4G1VZZq+IpR7
7lEaw0wjMAaojl4lUeYZxV5X0CycN8N0cBw9u60S6Mm53+I/YgJNgrs1o+suSFNYi709AQnT43Dv
vA9+p2mSA108oEULWhK2+kQjBOuWm/tOiSN1405gpJcxBj3Xwn7+ESEte2MRfsRKF6HmHqpjnR7k
B/L6IRGRmqQiR7r7SWMfWzTHChC6rUAcJKkuqfKHGCm7ZNdaAfR+DDmjYRzhabXIDPjyiYJC+daX
84kyeVZqZT3CJa5PWksEGwcCAtUXRtXYuf6dykqyIz9b2SCs0j4TX1vUCsSUT6LMWqwYAD9PwLp3
kVHbgPBvUVc1jcB29UYKG3t0KOX6nMVnLjdfUPBtKmjbtcB41UwBgeNMtKejihRhvDtRYE1grg2F
6DZ4tcP77BWfP/W7EfJuyehd8URDTpBFTDnsBG2gll8CNBwBndP2f3MaQoPJaoXVZz0jUWg+7FLt
K11hWJd6tnhK1SUT0rcEbbV7I3Ywdz7yCqigTcACmY0a31XyOpCaBLSUw2ftQbIxZt8Qei5c2ZWQ
JQNmXznCcS94X2DOWFKce5qFGshygB/R6/kqrvbJg0ZLWA/Go2ExTMaXUp1eFlp8saz8tShOW/kB
0EPaqIZ8aoY6cuJpgfM3WXS/S6kuBwxOSjivdbVcjlXbAaD0H2FIjInjohbrpIST1g/ASvqYhbSH
ClNSkdAGPDvWHLP4M+tbp6qt0R0NKolrD58EWvgCOaCgFkv2TeanpCLVAAbxMJbV7spZd2pdWN9N
KKZfwKEiqOB55xWraN/16ZH4heTI8philSvyMLQ45f7fF7uVDw6jH/6DwIQN6svpGxvGsOmHqZAN
gN5cDDQJNNyhrejZ+1sKv/5FZDYDDMBCHbSuwOxVokKHz1cXhi9VhHFPdYmLyCZymm9Oj84gIB8K
dixx6QnhqorLJnzO44ji0ZK83YK6tAfw5HHNBc6/s7i/BlnsThklPo5g7uwTQqBd+O7PMWtUVKOT
Ksopz77BSMZ/Rks21snLGQHeTV7pjqmWKEmVgilnmbJfTYjRNvFvgKXbbjFn0cPCl2y23MIC+rKz
cFaQT63Qa6ZmFhWyxsHLeMJYKmH4fJOmdMFoWUF5qbR8dSQj3wGNcrhSXZHbcpRbhY2b6u4Sfe7n
V1LrqC2q4PMJmsxh2oW//8CKS5whBLmqN7scYqf3foBfNob80hIJxMw3WzZiw6ZszvlVeHh+ZUVU
KMUsUP84Ots5d3cHGEOczHMDFCIA3ovdnT6GTX9M/4NSAj4VcAcQlKR6VP2SedZ2vuxIJvzGwmtk
uEEiFJ0DnsizHzo0drfJ2wn4Klkvsc43mqskAvBLa48cPj9BvejV4UWl3UYw5ANYSbZM0tGmRYXJ
6Ya0l5UG771bBe5mtEjmvrjGdnXpzbKRGeWP2HVeL/WcgWlHlEeJ8xbFX5LPszWH+S+esxr+Pi1/
m3tNLJAJVPycJvDgxVWZAcslZIgi+tjbE0LOQEW58J+wmUiOFXuXvns5NcrZn5dBS5F+zPIPO8Gy
m+TkSd18FG4q79YtODKOIoQaVT4Xe8YNTvhEZt+3tRdna41zGNUZWNzf1qy/nZkXVYDBLLzyT0+W
Ipt3F4VSw/5wGmzksL5CFeMv7hKXcKWI2atRFOK8E0MeCV/ASSna6nokcHtGva6z0GnvtUNG2+Dz
g+ghWZLBI03x0G3aGloYgFYSJbvpbGL67kyIHKkGgU3ajKS5UgvnDBYmal+tmL/4fMvyMo7ERzUu
2PA5e2xmjli4wHKK/i3B3xVKKqf89RDD+Gc6v6zK+vmVNEd8PLvwSVrVNPiWtW/+FBqTHJcde4rs
Ubwo9k5A39wrRXOlXdELgYtP4Zeb7WhBElqSb5ylVxUNHh9Kvx3RbL9kR8n6HxPGgCjZgAVCBT6r
ikVCM89ZTXaseE92bR+rvEuz5z929TGNk6VMPL5MFK2PSc/XWTqPAuu5xhNVjlUP5RORGzagmbyR
HFs5+JUeFQZPwYJoYwoL7sDqZgEUZLV4cVlofjH1lMU6H352CrFd0IdgnMXcj2uhcFENITv133aP
vV8kzfr8pW/Ayns1/ddsi4u3Zt6abMQ+gk8JvKfKNPpZJCX0cK8BKtJbXwnxNf3c+/m8jdgCyeRf
Lv81dYA6UBJuS6228ljQXva7cMKHFMfOuDdM7n3N91uMOQMlM46V2K2G6S+s6NE9XhAPbZDSXBhb
JlVVvy3EoO0Yil1hDPQIvIJxCgP0KsWjL6MClC2N/PyU7YUO5ZjcgoenDtKcEaQf36wjGr51Nt4w
9HESVxp1zvnfwlTgVYwFltSrG5ySjiLPH1+JrAg1dTVdpXBgktBSTl4Czaxvt7uzyMWy842Tw4yd
UHWcIEWiUIp4F2+yHYtZj25L8W2TMPbZ1QV1q1AS7Pil6w8CPURQCFDVs78GZTQx2pv4WBSgAhmC
9F4z2wA4cP22xYBfMBGaPoJLMFpMqGAspXq8DYU2g+ldJEsqgLBUaFY/oYe3wDBfaFGms9KkuEF9
IhrIIi2uIylVMGDZ5bA71kYT3j6Yh1OdfAxiB2Tiiq85vdwC5JcTdVKLfbanmLwsXIZMYeBNfgpE
NdV0mlLWjTgqOX0YqJwW0Vblbsxx0Ugm6X6EI2MRLU6mdBGbQ2xCW/MAcoHUdvCBjqtq3Eii+rlx
j5AwXvLR7uE4CWO0GZ/x1czEtmGDsFW2ohR5mN4i8onleRUdNdf8fz/Q9M98OkjoMG5iqGzIMMer
Mvus/NyKL24gmaUMiznOEDzkohcZ3oWXaaBbRto0I/yaGi6iA1AffJ4mRTmtDBGkZCXGmrjOefNG
TzTjsHkyveAO2DEukXjl/uPMUaTPND4QKPKou6T9axP/LLgSeJwnx3lQadrpqJdXBzgWX5oUKL/p
tPrFcam7H3GNWbPsk4Z3Z00EeMcLMTYstyNIJedebLEtMTshmM4JBn6mrfLQiNGfH0UYxvafbx0c
S3EN/e/N7HEn/tALNHvuXV0PjrD58haUAqxmzxc6YBih6507RSNRoY+0VwtFYiHpMnlJ1K4kTjC9
n3KhUYmH5fipQ6Dlvb2kh0PPTJwSuyCPljBiY8UuEYZZbZnNCPbXRhqwrQ4+pbj2tukRR2FE+1M4
GwbjobFGJJIAudlxV4E4D3WWCGQ6OYGUm/67iKUSVkz2XTe1M8R/gQCSB/qEn6sDRNwVcUXUl/er
xyCQynOzRogc0X2jEDIvOwyUOAx+6JQR41ZILzJl699DiKqCfzw00UApAsM+nFBZxvq8fMfU54z1
OjFW11eI73RMpP4IK5K4NJylW5le7N9jO2HA3uk6OxqG897qCX8/TbUDkfD2DgidddRRVIL9rJqm
juTNERu2tlVsDZxKeC4arEyASFgpAgEwee1YZCbX0eEcyKekbRXPiz8du9fs6uRsEDURAZd8oPiq
+MV4yWjBZzjJYfKghuOIfJU/lalJU7MNkeyg2QIwWlcaXiUVvi27YfNGhZRU2ZruqpwZsbSkvxUc
E/+pXYRMjK1W1U7a8py8CC6rw/4XGpyg2ABsZj99mTB6uuA6AtyIrvDEh1gsn7pyaq/OqGrRjNL6
uQ9mCoVbvwWzLW5JyKUS85zJW/NzXsxbqtFhDDQ+2tyT2HhLtcvGk/ro5mMlWY6q6ZDNIj4O3lCW
gIfugGMP7QPbGbSSir8vWkZfqwY2xeqE9yPoFolsZE8Goj6jrBSuyBju9PAxoZmN7V4FhunTfyTT
6wVKVA2zRdQdmh7OkKtau+qij9osNMUksxk7WoefZ+jBUyc30HeOSmzeW2re2850DNSrslLvy3eC
HMefbY1KYLaMQSu+rzWxy/LfnFEQOhZ4mfzXVUtZYwieg/QHCgXzaqJG3Hr9NIhiCr8VON0vldTO
1mg5NGOfsqIkNX5Fg7OszJWRnOlc14Ukx1+68N3zrQPkiuU1Zn/kSbEqm/Wiz0LB+AkW/861v/d+
NT5TcOtsi2DwI2V4wR9VBpUGVZZJjSf5qEY6AAK/b0rCbfmygTWGrNX5iwAxnx+KwBt2RtYdfBSh
kfiDa4QfCEj7FEDWHBvS2w3/TX8NFEtHy2pn01e8X0THMkPpzbon4leQSltAvT65QvsZUvpcQ7Cm
2mnFn+EnZisA3I25oq+ehVIV+RW6gejAQnlsMhtlPT3mdwRi6INr0BM4IWMPYy6uW34Aw+kgZPdh
494SrUC0kTxw9fZPN/+2jGo22bD4DN3Dq0zNz5yCGV27Ck3fdzvxC8+GBFYHp008ehI1WUKKO3RU
jPaoo9l7ngauZTP7JJO7zbIeedtmpqiL2+kuY5aoIVrlt8vfJinOwk4kw+FCSsmNDRsMasxax4YU
/sXHmio8R0Yonn3l44sYD9P4XQEbZhpbSaObWuVwqaUmimesIo0ph4lob2vQZkcB2v8rXn4Rs9Gi
sGKs6CHas3YRJP17xpbeFj8W4BdhLCKqWIFsD+yxtMCbcJIi2M6GEM67oAkXoIlTo1KDb08+8kLq
QzueF/i8bR7WlD91j77G2aQAZ6h66GB41J8EmbSolqzB7uenlKafiLxcPf1O/TlgqGOS7+6X28y7
VzHUHlQJ9ea1CD+vvHsDJVNhvEUHRniirDAntM92iFeL28FexIGNc0x2QK39Mn0H8YpNg37zIfJm
BKF1DWCeCdYxIUp8hFF3Zgp6IQ1KFDJhjVQ34cpvA+40AlTsJoHkMGlwXY8B+bt4mmZ6S9/hAR1d
bXo8/jLfke5C5/rJFedUar7izc+X2BUnoxbq+CY/P5EwniWj3ZYgp2TLAu71wv6kGGq8OTOCO6Al
NboJ/3mEP4De/6pNnxl5qmLz6+r+wU77NbdHsqdqrFRan8heGiwtWu1PQeqQpicmOCgFrnX8Y31T
NFek5VSUyeYzv8AroI3D7/q6vPmbmvxdBLXz6REJKTEVNRw/hKyyjg0ztUw+Wn4ZPUmAD9Az3W/e
RFQzJGNQx3iuCSb5bLTD3+htx7Jtet8bbm5yODLj1kk/x9Qi6Bg/0WDcwliHt9WqI2ZVJbm+/5XT
ZtmZTt9Xj5tu/MtsnC639aEnEXCE1WPDXdx+teemMmRWu78wwSVf48J3uXEXUk1yh1AcCQg0DDFR
utpnqWwHh2jcuvsOT8RhaJXAUIdkguQ0sWye1WKi/wZqjJ6wBy+9B+Kb6u+ScgUHqpvGtbawlg51
PviR05uL3K52BLU8GhWRFyKXR9JFUw/gcgrmALiEORrophGGNp/FWLZFA/AoavHxGltOmoBSNWfT
ksWAeI+jK0ey9Hx9Epb9RfZgZURU6Y9/j0Z0QL6ZCd5+vY9zLnN1M2gwH3qhNBvGRPFxvQZHNSSY
ukNoQ0O4388T0aWIRpC6YP0JZTtr6tJkxazXKtKvW6f6iitZc+oHv53e4XGzG73g3LAuhmUykSUk
WMDue8Oh237H/XGzJL56lmFukMMW/ze0TScil5huGycq+6DJHA6k6jqHGvjVA4+rnBnyu2tyunIF
dOo87vTx+I9paPPFfUgvQaHSHC8lGfiB909YwQ0e9HBORkZsEP+6HIdVqGiqs6Od6h+wY3x3Uu4n
iRK5ZhZkFE2Rh2bVBzOf/EWTo299+FDQnJmx9hL1617LCp/eoE3gW0gxp71JIbaotbdver1cu3Zw
I9uWCrQniKRV1Xy4ExooPkvpmjFZw7b3xeOM01l94L3CKc2NfIh0IucfGZz3gHueAai9IfFrd+Ws
eHOGhjRjjopQuLavKGTCZ9y/QE/TEnhtTTH3eF4N4M83MUaQbEYw+i8xouUgwi1Jxfus4pFj27SG
I0IjD+bxFuZxu3xQpccWcF+r1vFrRsaN5LFpTZlC1n5E5vj9AU9iN6cKFLN+1J35q014RXf/sVuZ
qpqtaV2lJm3V90jNZnvchp4BN9IkK52zcwXLMTTGVEQk+vKnbhV6Ei3cYMT7FngHD+kOI6JP6GcD
C1ik6P8mT73fHpINAWE84kB16/ZsfRZk9vxuieVyhQOWc3d2Nn1hDNKXpLx/wkfC36uo0Bd/ecBb
EJGmJB8K6ipy5XN7dNW7aXuJmTnr9YJH/q9FP5ruptU7YtM10WrsRjacP4e7KnyJ4N4UW0YqUOlu
yN3VB/bWku6KNQgoefUOGTPDp8jJ5T9/866QL8QcheBIwJBQqxwMtmkdhNUHJO4ggmXAL1xMjuFs
j9ishKP0/39qPoJ2AI8a15qE0pqmvTQlY6ejonOREwPaXsjMiQFDSJlapT88yBC3siTwfmyyFJD3
Pz4LTcIBMmGXPUzWAIEN7/tVq51VeuTPhyVtXaz8iqf53U39lYt4atr48EQbZYs1bVA1OZwAMrG0
LEoQFkkwp3H3WGuLjSpGpl94EI5fkoxQSzViLQtdd11QZmyOElJH1nGYfW6X9JTq0rEh5AaGsDrm
ReJ8eJHGyqQRoXgh65+n0yeuAeB4S9QBOYtbMZ8yxROmk4SF/GoZcg1jbkCBI246Wc3vXwSRDcSn
//nPGZ+BVCn8oC3L5yOQZHwWpwgOmYq2dYEyMAOoYn+qLtq1aZRBCGyHncuwlPiUYM++z0u7zasF
QoeFArX761NgIOtZAki7/GQhkLDwIoF7AQtgvrhfGuXTL4lC/Smb3oYj0iiPnhytyQVXieMT0KBL
J7e8wEP608+V/ZIJZULHAAcFx6Z4cyQFRlonadFDv+hVF0w5M07nG5WhJsZ1SUUnqlCE65o3ta3H
gpy5bXiPatHPNBo98mMegmuavjHehpbDskgL0khfmmZF+Im1FRxNWhzEe8GdkIbhdiONmQBDvySu
2QtxgB6fdnJDM1gladwqXE+jtmCEyMyYw3xw6y4hb7BNawQYE11ajZkZweiJdqN0wJSmXbaTo9Zm
UqLoekFCiuySNV6xsiN2ROhTrV5qZ1Y/Rm7l9rMK0V8DK3sewfvyiLxwYywH+DqH4lM8+AzitQl4
yZ2PdwmyyKz0wUm+keSI8Kv9VNuIeNAPmUpBDy7NdEHv0KcxPSSDupCdVUKvpIANp5bHxBjh29Oi
UXccy4YTCOhpIiZdGX/4L3innYx8hPchpl0LHGAcS1zckFqkYcE9IGM0PpQKuYaZGR7cqaCfcvB1
YkVZJo88PfcAlruY+hyste0EJOx8A+fQ0JsrUKG6O49E1lgSHXqr/Q8ZeWPG/kXp+hrqOoI6XLOX
fQZ5nsg0k56/8Z9Puib4Erk60LaxcO3w1r9hzkG7IhXomCBR+fbRoYRANDDTK17Wh7qsJqxQGu7Y
BanIRQHoCN9jWDzfmkMq/+zsPWkRZEEaPpg6prtewUdOyNDdlFvwyeZODUKl0OUVDlf0+ooIDMlP
d5ypQsPiDmlUUdU9/1RUBMTn+HCj0ZZyJe4uUHcUkpkP3wPOBt+kd/85uBUMFFCOyekczlGspd2n
1l85GOP/b47OU/r0wyYs4/ClpK0ZG5X5s1SndCNzrSELyBRxYlr2wMR9o/YaXc9j/8jBI1ZeYTgF
qn6SU2PTnKxT8tEt0EgOKUCz9yS0WC/URRRPpNCOuXS1NKx4bNbiSa9SPsVKEnnR/psTh6QWloC3
AO+WqtkU+W0zOOGmZODNFnV/cifzxRNcfuvSpBQrtK/IlViMmdo4opAYhgMyhabXnP1MFQ/njUWK
wyS2hiWyUcSka+dhReVjmIIM+0/stNpEB1X9XW4K0CQPx4DlezWNYlOhcFOqhtK1ju3CnzqxnXuD
nFKK1ZRHz8aL46yEgYPSIRIULOma4f4T3SZFdLHOFFrH8HJhBNhZGwnoQW7He0qQKoK0KuGnc3TY
ORCSDH2LNCg3MZVmO+L0bvkBg8fjyPodNjeQDSDdJ1X+aEFKOL337T4tY47sG5dwNdtUf9JOeDc1
Uqy2Mhb1XSOcxKglz+pzpTYECDqNth1Ny8LHR5hYlKeOFXwox96nptoQ5Jw9cNuk/5DDlxtgf0UM
96Hvm6dubGBKxcJnQ6at56estT/15QdFPPGhaO8IAZSaRVJJquV0r4G9Wm0WJ8Do9i76QtYs/qcs
JStkmRGTWtJq14DDjNXl7+Ge317p3yoiedTfPN+07R3LpZHlCUP8FZ8epS6WTNmxe4zhPkbJPiZj
9HiLeVBhndAuwoOvXhJq9JkSp9hK+/aS0/7sN7nRz7Rvz2roon5ZvO45TYZdFCcXLqGXFkzMnsD5
ZkOUEqRCJd+Ohe13ox0K7oFUD0Ry+w7HQcNxd8MuDjqeh2a9SactzDCzFmKgivmAjqxqmwl7eRZG
lvg4XBVfhxh/8EO3FB5zjplnugovl9jQ+IIERt+o22o74rUgn6wRVytiKjghJKy0VukKSP5baVXy
ao2qErt2EEKvrQtRzZBHdUwl6Xe7AixBC6qGHbh4joxsV7HmNatCD/s1+6pok1o/7Ef/QSwVkv8O
PiS46HJ/Gh1HMrBpk18uXSdfgXx0ke7TeBbACJzM87fU+UrD/oBw9ExiV4bHxJwyQbJOpXax4VWs
+NQcb7fiLxNCuNG0kmattk42hw3QFnfGxGOcHNiBEbnfAxdweb2TVi2dBAiERCRNzlnP9ft7ztSo
TTPJjaSQOPLZYl8v3FGZi5t3PZDdr0FCP7/y1n1JSFf7aM7S9enbzq68shZAF76Y+dVD9bJxbbJO
+4faemtAGQ0Ly01IhQVD2Q25dmpQyxyzf8e0dVpzY6xPjIaFFxA1V6MHvjErz+WqBTRlk9KOpZUU
QScd+BLA24luBzVcZ4IT+EkqemavcbiYoyzN/cldg0zGN3valhcCYMfIFaPHExXQtBGHy2BTJop+
UAIlLhyZNb6Dln2IMNCKdK0svVawrM3bKN869/zHomPq+Af70/az+dO/SxUc89QHl0f2MdJxbx1k
QXIlvdPdVwsL52Y/oqBhPO0+cYiF0VwimZ3p96wyowug9HKdtwoLCUF2s+8nVakoogSlUTPtJU5L
pNHBTT1oLJxhDbo9q7DSOuoQrsvLtHo+++6mVn7aIy/UwgCNHhlPBDVzJHc4bVNxHcXYBQjfSzJ6
Rkaib3REadknzEFXYDLCfF81EZK3SuqQYe+WS5hoZo4L/05MTqsVqif2+wtj03MjpqKO6yhi42R0
Bl6ldKqTFJUKqo/MQSrqmH5PrrJIqGoP2KGAM4CR2PA40x7DJa7aHVuBLEDSCwPZvKGIwtG1pZxc
973rQEKwKZy1mSTMGo6pgpx2niaGYajYIRc9dVNX4RyaSpWwkCGrxBef3fdG/NWIyCrk/wIfBcer
nSd2Pu/xRFhbwR449lq8oP5pBADuMRm84as/jQLArJa9e5IMFQXoB8ZIKciFjmob69R4gH2dtwJ2
wnsjYEEAmqg/6CjSjqIuid0BXd8HBAFNqjLoyNdkzXuM4j7Wj+Vkgcb886fSxpRK5M/hwsnVM2Pl
PNjbhTsrmYar3mmqZ3A2eraJYSaj/5uVKcHL6WSVY1g3T9BK+54RPUHNE/zSF8Ly1wYBcn5Y8Gnh
CBfLSvmtgv2uGzLsvpSnwliNFswOuWrj5uBo9JoUuA6WrHYm/F5sxWjwRWMNtpUY2h9ul6N4CJbH
Q3ua4L3nSi6aIuM2SonuqU4oHm2rjbfcgY4C8KBzR5t+SA7z8jJf+30AxLL51L+fC9eYQPk0eRaE
j1I0nXynRLDbTL/tcUn6YqFAHrW8riaBdatKsHitoTGr8GUATXgc7yRfGnbOSRQ2Rokt6GeP2GqJ
O/cpDFYGBxAz5jk6mqkK3S2zv3/f1dq/W4qnoXmX7AFVrmT5O/WeZQMyYMCJNDMkVf1ycMd9xL8m
SRSzjPu7+iIXg0PzYr/RgvxFouXpX03vGmDdEIxFImoF6XoyPTaEW9qqYvtciXL9qIWDQ17Cpdlk
NpaeZeWjj1nKohMIBidgZczc1amq8enqJzPLnbQXpRcTkMPwHMKtKttjJ5yIWD/vAO69CPyY1xF1
VTY3u16TR6n0h1oNocH6K7Pxf/CgHfdwMDhumaP6/DPLqqGwLOiAijfyyHU9G6QthiIs3bSPYMtc
WyxqtEfaI0fsDdlEPxuhXGB1HLfCzmxVELwAJx3FA4XxP73j1HrcweQPOVh0uOcKE3HzbPcrrMYG
K6DiaGertBZMRxRhgQ74iN42v6NG2f4FYEdtf/ZK6WqiCJibjv6A6lgnx3FQjzjiR1YBEmMV4uHL
XPPMIkE9uNVqUAROywTHWuR2Bjg1TsrUFZut28yOFV+fLBzuze60hbB/PdEiUbEsXWtyr5kzFYRr
hZLg8FuVEthwsyYRPZdtzDRmW4arik8Xl5oBa352AVPx3ZT6usLIKv91WW6Obh1y0Ie3qmJEARqB
B0p1jDZR7cRbVo6scfKk+rwzsVSZNL8XvH/1l/7ddfDn1CiIVApY0t6c32szu12copUZY5HCAXNc
LGxmI2hL5S59Sje79q5JuwZa/WRNpVW1SBDFhBf0VJP/tXN52xpg5OVWwE5uuMXbW9zU8F0DV/88
nnXRiqnNCMpYUYA0Z0lJfIUqEq14DDddzhC1Vja1YK8dgybyFaeODDUC+bYIsq0JAUSQSbMqkWhd
U3gKeCgQ0p7ynXpQlajX7oR/dlq4Q5fs2TQT147BpsotbTa1m3OoFdnxtpN7b3o+LqQBHHBdQgFH
zbacruoHSHHEOvmeKgbSyrDxiDTYDpOxmerVOwUY5sFvqBuKEOh/4CDnEA9j7FFQTcWly1fXPKEz
Z4u8cf5bZYejIrAWXuCQwk+3152/5tteW+LpmWrjhpUobYseDf2rYsl7WLAjccy5G9g4b69L/v+H
Ejxum7M0L7n9RwoUFEUk946bFvNAY+Bg+ZtSGKc+im3M0YWX0fhlbhmNncIySH1axiQssN7Fx9+e
ETlfApz/k0FYz6uPDLzuU+2Xl1cyH3YdFLYaUFmHYkyNXCdjq49RKSAod1CtbMLDjChuWq70r3l9
IYFzEQfVGl2I4/xdgIBee/aT/qSg6712rmuGx2aGL3KRy298aM8L+1J6Wuw+FhQlYJslJAgF40ww
QnoJT1Jo7seK+WmWHKa2NqNGV+bxXd+m95R9n3R4Vrg7gT6OJIMbFfdw7QLG9FKXkYosZEKBd/NM
ClmNba6J52xsPj/vXl7eOjjEH/iLyyGxcdqtm9zLpKv/BB3cbFamAebw/kC7E2BEt9p6z7fEW0g5
yYsduHrAUFnYlSSgHmGm2T9rdFDBBkmpoWhTn563KOfMT1MwEZir0DzQGO6sqTPZqmAHrLVDYJ0+
mbK+KBXOoCKQixpY0nqjyrWinkGL9AgQSHvjAUxVRO9pAwhe+vOc6Jmo+VqhjI+uXp473Q0f8AZp
9eq5ee6wXBM7BkTTJ98F5T5yp1KQS2u5vO9uWlgsuVwQzWLyDOrZyCqFgO5KQ7AqKQ0ADynAX7B9
KysCErvODZ0EcF3JjIx49h3rLuh8pNFzhqsEe0pSdwdJ/OxxfnuzxUyghepD/y23++F6O0JlK1OI
Hz1hxFE6LA+PfXwqYDLu0OYT7yQHfprARISmb9qQQmvpF+lFEqVR8AWwlNK4bZ2v/I2Cl1TK8PAl
pamaDRicX6f1HOKqy2NsRE7qTJ0f3mgfhHhcQQuYfjQpBSlp17OtYZI7W3ibDZwxNrlZ8utaOEQY
jWpOYan29zxuGIRzM9UXo6hNJPswHzIhyEF0TzKAbAlYUkPAKtv8bGv0ILzmKMT6gpZqOSz8IHSP
px0Iiy1gcaxv7QFXKprv86jcQ1yYWBfYTY3M+F8Grv2qIoy9nUkL6dNBFin0+UEMbIggo6R0v1rN
5uqo8/orTNlRgvzZJJvmUyfZ07dcMHf7f4nUIQoZzmQkZPYx7KBLR8o4piIVEV5U5HsXYyz5XNos
oBBg6OVLPCTEiZMwoQoOYFQqmFQ2vk4AVTTaqud8hg6YQLlmCwdvvfMGSLD1zq5U2yRlRErjwI2K
kXu3GlHpq3z2uFH7UI7rTkCtl63jWV/YpTicUyw2XkB3ZQvQcYw4Jiah/WSZs2BUJ0C0WtNJ2VYz
w080FiBCOtapmpp50E+FEoQEyBZqpLlLQhyIcUNkjaVIJGbp9RdqmNfM6Ol56KkVO8iDC4cIZLep
kPbTL/S7V525oatg6PtYdSdocWHvgh+fdAf7uY4fOH5uAqynhI4D5Y3HqmsArF5b3kWW5fYAoUP8
Ma7bIR/AltbsCnS04hgSmg9FaTV7/u4Au5N0f+ixuILmJppLZOJ6D9CDLWdMnx5D4MXdx65adnx8
Ccwpgms2XbGsGMFuvjn4JAz3obrycohj0QczDhkFdde2VEm/3JzbDqf4imvmSZbevd2Vw25z8cs6
KBoGv7q9IgZYKHsd1Xj0I5Er46sEW+MLXZyk4CRBKF6PWiLVkx0viln1RpD549m74Dl1y8kLDTsJ
IkUs76scrayhvjYnUO43X+XicipPa9BwKmgZtpguym/sVXWo4UtAiFkoAT+A5OMvKLVSEdRyMc88
pEYUcWFSdoTF1XOKxVR8wXwpttLMBJw/tXA+IN2x2MFevff4rVhdQfwstc1a+jCJlMhL3hY66Khw
x+Ix/YHL+O9KatY5OTA32tktYxCC+TjTe1xGBvT5bt2hH9ooZ4DLOPiGg2ZfRj91b6mgDoE0bPFP
GWxg1L1kjuuqUrPNPwVrB1Q1MvA3VexhgaUrO8H+5vktvD46dfsghXsjR/HQvnPGfyJi3Q+n0thl
RF1jKJaf83Ha4wq6IZABbmxurpR6sjEWxlgBAMhbjAhEfNAeHwXF7N+rJuh4NRksgF9jbkgz6q2p
33a8U75hfJHz8RZCmnWYDCN1DyH2VougtHbjQzc+Xbzr16zCXNGm9cwPEea3pH5WkoNxASqybgIp
74BNOdss4ghWbeL4oqr6LVNBuCrX5cDa1mRsavPxhfOSOHn3Zi5+sqsgKXFcCE+qL91leh31aAu+
X/kGpiw+8i6CMV/8gRn5Bc/YWys+oyEcIlmzlPJF4Ke3oozofFC0oK7B9vUfG8E8OeVz/AFvTfJ1
o8VurdobMaaBujSSG2/taF6hNpmdTCCHwiNQFP5aGsYx8PyQo2FrDIfosyuXDEQdkox6s0EdFMBP
wWA1tOoyhI/GzCcIs5RtnjCP+ih5u/YA7sEeoSLB9Viv4iWvUkXyUtZWcp3HIPreShaLz9CGbQMc
km4nf9Mc3f1Bzp/P9cFo2dRTtYZQIlmKLuuQn+81F8YXR5OYy/RYKHmFNk58QfLWaXF4Yo1hn8TS
Vhyxb2Qb3+81oZ6RWH7e0CyqB+B1lSlhQPDhZivsPWJhMi/pNzm6DPSw97CXOuoI/zdZaYFKhciH
LBuTuJErwwWWGNZqR7usKZzWp9aDpeP/o36gNvcsJfqXcHxiz8qcJpBW/S6EkWjlvhYw2vrz3lzv
aSaUSbEixtfumcCnt4MEEpwKDkwtUdkbWiJqYNjaaak0ieu6YwcT5pMK8LyUHwgFUnsvXeq9MpI/
LJS8Bi3Bf8rTyj6FATEGm4pr3OqnSFCnTe3EvpeA0ZHWxnIzT5W/R4/gtPshEVPhFTnoZ4yUSjwq
A2kX4FWxe93CNh9fWzMK5KDniUrdE7LpTtQwF1ETF6cuIxO8yamQ1QbIw8AOMTyQ+qqVggiJnARE
Kj2jR1qHcfao3dNsxwlrujZwA1I+uiuTWygldBqq1k2uVAL1JBE4vbetcTq9LCQ9GP4zh2AZiubM
8FsFm9DsDm+j/yPmdNmB7RPVZc7gz3ZsSAdwYoE24OoXqixEf9GazSWDRwqKYtH4pIO/CYAnpUFZ
rF5RG6h2dLhBXD+QLlhiKYpOmerrhjNfYzvMJP7N4K+q3ugOjJc1am+kS0JUtgzSl4AEK8vXz2OZ
K23Xn297Hn89/zIn0dU/DLcidagDt0h8jeHM08jmlyDlOT8tl1YVqGrYNG//FOH88dUVN436B1ea
9Cb7Wj4RkQewcMP1JoArwCIZTNa9oTi4rfaPdRGNdWpukPW+Tq/QMXp81HHGqWbihNoYLHdt8HQ5
neyV7cRK4kidtEUzhRH1wV2IBH4i5jrC/gBuPySfTNc/8vH55pa40LrTqKlBKUzLtiYUBrEVA/CG
HfPPscOqWZz9jw8oMkS3izLjqxYdEWSYCZboPZddi2nhAwyK58jQzjJObXvZHj142rgKW0U7yHWd
lGekK+C68endbWN3hitadIangvVcmMwNrf/8xpty8gCzHdDJ16lZxyaGQSlq6EKom66Hbj3dbDmJ
ZeJazo45DIvz7oG4nd58oFLpXZJajtAoNRFkAO1to5Wfqg4zbDSSOohlwSJqZnW8D2Iatn3RYWy0
BVaBwpmP4ZT7+zs+FvHHAyB87/adDXA8fHuYXmlXL9BsbR5Y7ewQch4BraZmbFKsOp7N0SNrKMnw
eKnMDSLckMi1pV864nsFgx6zBWupoXzZRb4vJT4jcDGMlgMIJVr+vt/J95z8VBMRFe2E3t6tMyXk
iFe5Ca6eVA/AmtEdWnK2F2rwAdkQQAV9ruEsxWST3fi+LHt7pv8im76T4nokZO+5zlYUm1Vs5iPQ
5QmakwjNeqdmdzashgsAV3MgRv3Pfn7TFGhIq/Byr7FdYG4jTzSYMImiSYU28T22kHe+JBuCTYRo
UE/qcBmBFa1MPks5FB4ZFB2iN91uTNxs27Kg5arU6JxK9T6KTYxyMp+WLb0Dj65ikYVuLWOFCP4/
3vhWQSo+n/J/ljK7/haA0ev9wMwpFkR9WT0TYGhwDq8CpC+d4QYkyNtqxyx9G0i8baBXvNFi/cmJ
4R4IDIjVo5/cWTfwEd+cMo6T4+DM/iDtgj9qmQOT9GBdCNu4btZlNRkoWQ5KbVHqFF6V6+GgJr9Z
Ig6pxIQo8R/i2RT1icQ5U9JBt99mP2CVzLphI3niMQwILCm08OdJUUk1DLCcVj+5nwQ7/4pThmtx
Eo+mHeqyGzcRmZLekgICc+n6ry0tio0TxRhaGFxujxend2mNoDrod/pUyIWYqw73K0ofchSzMHLW
jHWjvBnK31qCqeL7OcyQ2X8IjpOWSHf41wDJGVsP7YVyNI0rnpgh6azJ9wXGJHgcWUVGzXQD58RJ
sDAM260hhrdCcdYAk1LmhiHWw3bH26yoMMoeVfTSHXQgimfgsF4ZGfCkPglwPCrr86tWyLJ/cP9C
iPFXs6JCTV9HVuvLzMqHoXr04NgRYVCAyUKT+IsnxxNcsyY6s9MXbyjXCGbqFj0Ynsnh0Me7hsDv
CBBjQERDco5p86chlpS27SJIkW1J2FjO8SOz2NAhKMF3qnmmXMtRqvemzelJDerlAJxdb1s6LKJF
6QK8R+ODr3RznsaeGKISpeNQA7xto15B2BRhCmusD0wpbAYklOQdGWbJq7V4FM8Fe2xrNvY7r064
DAjXfeme/s98+cMZIfZvpQmLtQJP2Zi4n59l9QN+84JbJoGUxbpxlE5cR/eO04HS6dPoPgc5adOS
KafO9glR4wv+COGLjJnH+tBgAzR8cYRhhn8txQGte1+Kdda/ECYGKpjiOLu4vl07ZOwWEn0SgzDW
001RJsz/+aLFujQNib3QJNfLbMLQIpB8+YmiO3okxY/9NV7PEQrkAfzgR21YxzEGA4HyJepAyZUE
DMtGM5TV8aZ2FdACOmBrGryk58/DZ+SIO3QCS0hkGPiqsdaAbnHsk7sJlgivY0Uv5o5bfqmkyypZ
nnOUfUeyKS8P8MDOikpNfq8mlvqwZYkk6OogQbGA5XsWXKrLQHS1Rg+OUnU8gxtS28zmSyho6MtW
gT0+BD42DFOSbg8EDYD5b0NnIcRc1D2edQXWguivImm+jAShbr9CulhMk1OMt7EiAK5gY5HaQMDz
H//uB6l1iN/GPDv+qqzxG655/eB2dSjY4zSX2yU1NAVXSL49HDUGxb2z5xjkzEjT6pelSQaPAwyo
j0IQBbCdH5VjeFcmjBF6BOmkLuP6BBpXG37ES+Dya1RCmgZYDrJPKW2B3rSflJOmNHBxJKQrXcBM
2TGxrKp3EBEBXTbZXGWusGjJnJOXiBIcggc7kfaVJbgm0aToRT85v5G9oPaXggrLtmP0mGHHFOES
/COC9UKcNfPqSLB5jhYCHPMJpy96tjMu/HVJALB17yAjV5YIlZGdr9nxu0K0FJ6NdmaLUKo3s3M5
H0a9cv399dCO+69oKVo/1bbmO/0nh8Cgm6dO+sFVoP7OMoalLMgcb0IsBOB0NvX4RzYk9jWZT8a3
lOuI1tA8BScdupjCi7gprCEcaS+dtLLhvcbYE1jsuzVxCKCmPX288mAKcKPK4v/cCLuP3+XuOF//
XiNmNRmmIE+xfrBtTqUFU3roJdpBMc+aJ4aoZtBw+roClTIlmyCstVRof/Zv4BWpAPRif8qcSrBc
yNjdRMOmjEzj29tpkG389EGn9N5HCi7zkgtjJKEqP/rU4S3nwpp7mh3lmtjYz9Ifz+fZg8MPPerY
Re5P8//dDayFjvoYjQ7TnCLa6aLmO3s0KOlUfokJ6HNaxZCVxEERScHVpXfJbDE0yl125wZOdh3y
+tO8k9dIBmJIloJ1k7ITEznHHwJPWRmPiJZc0glqQ6Xlyd4O4/JQCO8otrAXT2sEftQTpfUHecCj
/TY7aUumXnxccKy8rFH8CyOhjr957ODcVAi0xTFIJZu1enZHVDs5tOoe0eGT3Jp/RsYIp0OyAp/U
PaQgt7b7c2nSxO70idFL6QmswgmbSPbCu3EKDUgKhOQGgslMQHXeSDKCzdiIs9dWKUgEvS00jN/J
SnrqpQZW56rR+1qmgBDNJsglpR6yyV5p2/b53aMnGrH55RN0aM/UKyst79ZMf7xx5KT5P3Oc3If/
mNWhUnTlTDlB0BBC7xoCa6N0Fs/7b2N30kI75kotEB0En5uwXRsKvcpgxhYZ5sb7sLj+hWvJrZ7K
1zyXVMRH/XHQFy2/EyzEjlQPXJQiJjpRjO/UTHBnwwM1gY+26PzASc6f7sZMcH/bPfvxRuWoCJt/
njRIzPvo/hvN+V6HENfIR5zSEH8GhUKOF3ecoHegMG+Kt2zgaJxRCISGNIsDFjUeexpCDs3sEy2c
kPLInupFWLrqRkXFwEulp6qryhm7hg8fogQhxlnmI+fjXY7eRto70rjiPfbH1CcqRObOD9qkl4b7
EgZQmjFvY3yg8BsdHMNP4KNY5M2oH24NsA2eRxPpo8m7EPDEgV6AZFXTsDr6DDKhAmhDRc80R+BT
GikSPrK4BcrLg5MJQ4TLdKAJM9aanHOXokv9mnI/5QRfUf7DYFxAJvjXqjkLr65HG4rqVfcAdeV0
le5kDxc9Ke8vBOf31gBWHtoE8JowaNMIYGc4s7gTd+bWBPVpUFX/oyNRvRRVD1wFA/biIKUJuA1w
Vmk60D52tJcV/OfpzV/Z86gEt2IR/JR1DQ1eNlWEJLxS1aZPcMkTlOPUBPUsIMK8kj3lR/Q64L6O
1RFVOoAK7HLRKt6O1Grb1AKWl0CD1ekKNoI3AGkNIq+l9qKszurhnfTBq1E3PalgPxG4XMa57BBZ
rrf/aOZ51WRyPxe+8rD/opMScZ5b/ONSN2giiaVm6tp/H3Rfx4QiTFLtNznl+Ok7ZChjJByp0sho
hbos/+k3tdLwjVY0QCWRVC2nyB8B6Ver1jCG2BMPVZ6+HDM54q3pWm2l1U8LK1CrH0LpUEsAn9EL
mcOOfI/b0IeWN/pF0WF6+g3JSTzwRRG47EvBQbacoURjg2oADGaccMwIguSNUnRBGcZYY7Zi6I0v
5Aj8liERQjtedzi34Av0EUJKLgQP28RS5Ci1hQsZhBRmNHxBm7PxF+xQmX8XTxrCwtFxvPtb6zib
W7tXhVUTrDa9V9JOhhYgJEqIhz3FFX5tuN9eaOl83cIvXgudR2wqEDTnkmxXyiKrKDNmflo1QZWo
1XP92ThxwvbQhCK2wSvsKxhC1Gs38Y7+7UzLapaaM/BVLaDPBBalkA23VmjHArwiLhh1A0v5HVAv
wI3bA7tPaIDlYtBd9OAB3a106NQXzRQ5D2rXcpnX6UZvGASZaMsX7xLNVA1X/qp1jU/WoHRBb7w+
fkxNjkiEQ18OGL2i84tw2zTP7iMKRXSQlQwR1tYVQbVQmbgtRvijem87zewq4IwF1cS2a2axrjJq
j2gB3TGenSOXo3pOgfXv8aNDsTUDYX6t0u4xqFZD0CXKpVRGrh81iNluN9Fl5YEeesWHcewbwNMl
d1FaBrPKljw+eU+kXQvV7H2e3ryed77xzS9Cpu0RPudE/EMp54TRMzsQY8k4l5+mXNIo8osqj7jo
d4DXSIwgG/SdW4Ee/ShwX/0GApIsr/fcAuASskSHHDI7cSofEoOBA6JdNwKDAD9N9eezaIkOXC7o
bjBRSERT9085Py2N4vMEK0578lZUbTaiQqtMbCdrh2TytSVYyZpbxmZBd9708k/U4YpvCzWsqmes
YHerXjJtxyU0+y0wAnqIFoiIhNdHwsGKZLTgTuTYlqrIZRHcTV/7ODy4UaFJ3ndHgn4W5yoNc2hA
ru/mxXwcUid6yXc5rTz/MOjpr0VhsluUWHhj4W+bPz+WUgS1n6o1VM7mhKVinCVGuys6KScdc7r1
i+dP7lMuBJSw9mGCXWs4A7PB7MdaO2QyL6oqCW45c0YsPZZHgiFQTdFtvZjPjskmy5anHELMw4Be
QCSV74rQtELG6vzKvSf4qTDBojYDLWz0faomKTFahJd9E07x5pdRl02EGqUc7J13OU/sDVL4px+r
HjrtQt+6NU2E+Xi9mvLi6UCG4jICkTzDqK+GIrYOQjgQ5i2cTaMyNIN0rOQemMENHr56q5TbdCKs
MQwlWONR2UI5bkA+WDFR5MCteXrZoqqzi9UZb0oOr0XB4Ki7+TXcwLUOyOAePOUi6JZy3nYLcFj2
3Q0Ah5ixT+x91/nsxNplGic0Ok7saNDLp/New55n68/0L8g1+XKbxKUawyjH9VRXRcZ3ykfV5TmP
9B8P4cb1HWPCf4h+lBSIc8ymvi12U5x/X2F6AeZGP+X5ynXeVJmbg+CWNsrNrgVpIXMTq6OpIIkN
4wvaQqzfL+Ft1G/Zfe+f4BnvlrKID/rwHhFYedH9Ai3aTpIAeCNHexcfcsJeVpulLk1GRE1K5TOf
rTuq09D+Hx/c9MUCHxX1OFjn07PgmraZethpZnQiHmzLTnWFbsNk7asC1XZWUE+hsi/ycXZNKmvL
X9RIfN8PhaFG/C9bgtsxcOPIvCdbuAmif9eHTeIX8aFjlofQWyiOqtjBr0eoG/fDGRQ4Y6CBt4BF
4HByFBCqpONnj+BUVWPT6ZRVHfjoy6vXVMT4W3U/4eYifI4rsP/Epuopj4Xn+jiUSeIF+ymYK3E4
VL51VALp5+jyNGK39rzPS8xI+3JjhIPk19lWOiiEfkCx8xP8sO2c2zXjtCg0EnYpSp6Nu7XGE5YD
z8D6xqkMUa+cEIakjlGWg/6MiSvTD7CkrBwMsewvJIS51zBXhBkPxQxVYmcj7d52POEdVQDkkD/A
90t2lybm0dQ+GESJ483bD5EGlRSzGAmlXQ00y5zASCGEO2Zj6lUotcY24Z3G4ySF2FGkUKwBnRgN
9D7nzH+8TCKm8EenrABr6OkpOmBXOfKpDaCdWJcsPLqMpiL40t1ASaui7dCokBzxDE4+6SagOUPQ
QSHnFEvLAGcmfvLCBui1fg+CB5YJzI9c+igSMpoE5MniyfMxXCmUscmP9Fh8caeQZI+2MW+/HWBi
OIGH1xhS4sbCQ/7WoCrixmGX3azTkGjTZOTQryy+SAcNl6geKCXQ6R58JpIV8ARG4MulrCFfv3kg
XVyhBIFRzpcb68c0UgYvz75t8ZH8pLcaykTaCuBRGpZtaso/W9d0TREUeyBbJDJXrJqj7pLRwRyc
gAc4s0ZzQdWXSSQZqHYEr8WQufzl65HcnjVXUbx3Wh1yhVdtqr++8osLF/telegk2+/+wYro071+
6NgyLryeerRQlI2uLsQ83OJrxTn+Ohq97gdaOjbJ8YA3YY9vawgOq5W2EkUa5a1zhZP0ugMoAlwr
dNperAf32i42CdpUq0psGr4sETjyKsKnjhLsZtQoNEtJLo+oH54RaVlmYjTptz0B8TLd0dzIX7Zm
DgMoufplZTjn7nBu105aEIVddC/9QJaXI0Zg5BgjbtywJSB7nWOTSqf/pWfWprQ30mNgDL1ASbei
axFke76H+WU/DfPbetuUMKPFXNuyj+7XHGBWn/MhoEBnGYW9tcDnnr1vllsUaou7v9wFYgrGc8Uo
7s04nfJDc1YZRtYAZB3R50weIEvPB4O98vQOG9HeX2HTvePItJUBo/QKHyq/22WG9B2UbQrPAxER
xq5GCFawLKafHNvoFJ/CdL/ZeRI06sIKjgzzHTCxwYm40RuJqWUs+6XT3XvfGjb1rKafyMeXw7Hg
1QN6UOe3F0IU8W7QnC1rAbOXzD/fj270mEt6jBWr1KhJq8dh5HF1FiRrCruUoCVgKPVZBg+RxSZu
ZuY1EeGtohRUgwebzQHeTH/hdrEDzkTuguo86a3IO4PMvCkudNxNzr2+VvRlA9ueUA8AtliWvl0a
SkGwlTXs4z94riI7nOcZe+3i76zdvFIEEiygxtmN8dosdFRVhGXKPn3QCTtKJIltE4/MqOzLcLop
nN65RyOHHOlizLr3fnhxY3PjxIpQ71UGNV+Kpti/+oNr6+ONwn4SdUaf+EeS/pR0Txy/mwVHeJmN
4PhFvC+mffo1unz/OazQZ8HEi0Bt2C7/p0FkdE7/+RT3o4i69M1C/o7sVUoGGINJXWlJQVs6NOm+
MU1twyPLksNX2NvzdZbvntOE6ci7BfP+lWGqtqq0HdOMN7tskrCCDVWrdFX2zLk6LhrbQ63zXG9i
26PxXJSbXgsCTS+yU1hlrZUTu1aLVnaINfQTVMCzXE/N72+9tQ4kpPdcx2WTfku7u6Vk52Mp+D0m
DE1yCA1vaj3vhqaAXjlVVkk/z9DWVCMiBdFQynr8Xe9N5JOtoJTvRJLI6Dn9WTQxH3Rbk2yt8tno
TMkufX05g+s4QsvsjO+lVcmH5UDcVsrPO0qUHQvTkCpsZyM3yuWRjqeH2SHO6y/Fj3PBmahKVRBx
dTHSZeEC+dZnXJAkfXCRBE/5ABn5QoL08vmtSGzeF92OEy4gd2pxaeXCEPfmeg3fPWSq9xvl8sjW
PCbZ6TR4EZ6Zbol+gv2vNJZSn2WWL9LwBrnX7ngg5zQitvqD9WnYXH38rDIL8vMfJi50WmVsYxhR
zBLyMkIxWIIAOZgtyOFWGDTAgxtBmBb81LH5CoUy/acOcQq8rprEsKVOufXW62GPzXiKMrFKlVuj
cpkFJQR//msCAUPGKgVYsa/1hO0F7+W+6pTxvojhCNB6lisyTEQfv8yPe9cLL5rjUn1l81CJPvFq
S0hgcGhVpisRv41XBJ18HxMDGG82LwhQmKXumrU/PqBQX/IWxJJmsEmNvgFfOVZmOSrGaAaZCXdk
Cb4imggKPRaNah5dxqOuwZqIFUsN4w/fAc0PysHnjTmKzB8pAe/pToa9xJWQ06QWEv9pbF85RPd/
+HyBAHMH3jzg0pJWSOWMg+5WlzPHtVgMwGMO8dQIpNrgHiU+YNGpGcvRSjJl2lnX+1OhTjqZieUB
FCxN/Nubcd9wIeyBdUAWCvIfY7BzVIjYM0aCEFa38yfSiRmBUDz4MEXyANOyWpEfvcXrPGX/F0fH
Fjb3TNnwejhkw3wWM8RkpyIh/Xkjar3uA84BQ0UeJaL7JAPTCko4xcGN84eWzsZJx65JH1Dp8xwy
fU5KGTeX3P88n3PRW3b5HD0QvgFQZ3889QODYRv8CxuP9X18coXRFiyXfRusAnekybebWJROmf8s
hEJbtM/7+miv9cxs/l8UhChUK/ahvj1Ht4C5DeymBeozww9UvKIywPY3N0fGvYlBsNiiZIU4j3MJ
QcrEP368ma+ltNBjYsEoyuzQDelj6cgLa6ECGJLK5yBkX9E7qzASQJ5+pfdSS5QoOZAu1jNSc5mc
3PQgBChKSn7oBodbv+2CcUKaUkY2UEWHS54klDJC0jud9ZXo9pO03K7da/WGwflmZIGIRWVGzwQm
/g+Josb2RaQPR8ctppcgshAlOtjY19ELdq+cjwktLb6oabImE60IsWAV+jyMkZsRpH90IMUgUb4Q
T3LB6BVQJ65/XBefmsHvlyjZbH0S1LLasmCD/XDDgVT4j4ZC20PExduiRQDsQnB7VOwLECRwipD1
v0HllZ97KHjxwOE9XBleNy8IDeIX42SQQJMr29P+hWLPQTIZ9IjzJki3CMJfcW7bKXDQdwQz41ww
hsG/6IZ0uzZ1T8eT0TwcUQuq4BS2szPtLZ9t7pMZQKPXUDYMOWiy377NFWb24UyDg/CzFKDT2WFn
IQzFW35dYOF0MZwNIYo89qsU5Hzxx83haZSL+ciBsMw4C3rXCm+Y0tJTQEPv0O/HRij1DpZUSWjC
HsiQNcet6i93QzRtQ97WgON24pMqlajAaE2ZXGbUp0iyOc2eiDjSQQQuc3q45nt3rDSjLfQK2gei
NWOClqehQqNnd56cBeZBpUGzbtMC4fca0jEUxMTkNbfjUpASUsxdIgFd2BN5DcCD/Ga76s6D0jcI
zTH+RPALk8EI3rNLhy1ztm46MZ3UA/WU3O5W0MPVf2kn/tKwXXJlYj3x4OmgTB1SXfskFt9LMR/A
ic6FGNHPDu+BARidhimqmRtYxCDXKnLcHaHeFeKGhYEwbi/rGvbKqU2K6t5u2Ngf7nHwIR070qZD
rXaNhUDai8rjzWEZvT4lIpsfE+nAWiEtt7NgxS3I3nRuDykK5TBfEAqfaA/rF+CA93RkAgaDijo+
on6eZtum6b5Z5Ac8Dr1HGBhDXqmKzoKVrEAsXhQAWD6BmsNFHN+PhbxhwSLovXtXHUp4T7vhh1EN
XNMPVHldfKiEPFOiUb7bDPg+bpWy9k9UpQe+Y9XHnSeH70utulSdp9AQKY0OH0CgYl/Zis5wNGpK
SfBH+u+ckD7nEDZMELnyPzbSYPb3udQO85/tNyHntSC6ipqbFA05tteZRY6bDdYHalJnBVR1fNwo
dQvfiRoB12lVtafQNaTIItwX6O5O1nGQWt22aXI/ua8ylHwAcRrISJvHctSmCCPIhzzzEo6Te8Wd
8l5quO4/9iQ6c6pyG7sJ/q6HF8jSNEZk8xRybdt7M6GZErlOsKiCdoO3ACO64z3D9KtIEfneNhkV
Rc0uNLyRszXO2mSMf2f1pzBbUoBXW6Q+5eNukkkfXnkRQ7H2N1u0i7f2l+8sRp/k6RjXriYiTw70
9y+uQc85Bi93b7OsG3/LSZIax+q8WR4uv5OtU2xZa8D3vTBYajHNzs1VbmBWb1eNFUfrLateya6S
cG6Y7zy6Oo3y3q3KOfawhEarWGOj4I2IPS0/1WskB4ig3N8Big95b+eMQD9LGwXdKcawo7o/RQZX
T40hl3/i+U7gUKGB+9uZikYaPmV4Z+OyaOBRssRj7azzOcm/1QmkX19bcKerkcfq+FmlNmeVyKD9
KxIhE3KYdKm5IfB9WtBSKWuDnopfUtU9Wo76NcX9kOU6RJylNZ9q8JrA2iYwHixz2jc4W1DTZaA2
MW/5U3kzk7PwRd4pBDrPu7x2FvIouPbwXSIg4BJyWAAVXjY9+tCkC0gHMgt83Fg8j9rQfdnBqFmw
/Uir/323O0biWdPxRgIeEa+waFR/5qfVGZ0RDafImmam+EAK0Few0eTnw1TEVQ0VLTyb0lD33iTq
F3qQrVHwMpOb1ofVTszQkXOR+6vGA3x7clIAqP8hMAztzjNdn/JKh8JHMobW8qF6x8j9SO62UXEM
6zaKqcbV7OrJpGTjRrWicJrnmrPE0WSJy/rXO3QaKMeq5Xv8XHy87a0yNpGYC1GX44l5EFqlRG+R
Vb3H3jC6ej2w2K67A5CAWlwK6YcAQEJ7s+HFBBzupUY1BJrxXsntXAIrcCly/CAeZi7Ric6T3Avx
KU/45IarX5p3tMu4nIVPU4Mcb50qteZPmKcx+9C76NiAoYa7uujyrwnMnyGyNMBph10qUvdvDEPT
IktZpkQTDpfi+dSXeVnUJIntnnFs5US9F2QPTrQFP4LalQud/0G5NsDql4hqdxeRHulUhlbEP7px
SogShPCvfJ5SE5NaYv8aKYOak8WEaohzSvsswts3WTvGsASrRHsU/f3YOnr9BjkdJJbxGapAnBsE
wK1dLodwvhkW/osV0Tt33QhIWj0xzpNdTlJmbwZ9Vnuf4UqcemaO6CQUyCjqNyFYZXKCDOs7wI0r
VxYa07FHgdIc1VDY9MMBJUToBF+QpbIjQEgLUgI6uyPwhVaau5AR1H5/k3NZqp0pZMAju6AIcqPX
qE3TxJryGPV69Vts+sPde44lY+UEtzFvnc1bHgv7lelJRJuax9zYmz27ezQIFg65MlLfK4/QHaeC
J0K0KOi1mjwRiJ/hGJSDO/r7ZUNLTMpclkz/I25RjjPjWs17KnNj+kkWFZuZTh+dPpnMNwMu9JcK
ducmn8lA6inmilKO2+pQFpi7JkObvH5stk8yqDm20cbm+o1FSX/0n5sXJ25MSyjAi20e7CElYNUk
AQvzkCclyLD658OWO8Wj7E77y9uF8xNCB44xLgW8xy5BS+CscyX1PZvUgmwHS9TKOgzhIstzYb7Q
W3uRBz7vXuf0dYm3VCfLD51NGdKyVYdqZ0wsyV0zU12JEEYuI+1WPIn/GeandJgXR1e6iBb38YkQ
tUxFI3gNL5bIlIm410rz0xWcwoYAT1v9bssh46UiLEUrxha9d258M00k7HWDm4PUtuf/vJilVnzw
VCBRPTPb/3nT9lge/YfnWftLnW//W9An7R0GSBu5a8nJWw7Z+tKz23cZRc92zwT3e899a/04avKZ
lR7rq+ba0ZlQw8rhTCzqKBcvvkOuoctFd3Wt2zV0ihLM2Mw4xXdGch3mRctB90AI81P7QtdxJvyS
zYt8pDdhj3ySuyRh9/Y+SKY9o4tO9gOsKyAHbBLRvd+TJmfzTM5QjKReJtKf1fbCBl4Bxr0gnuUB
3KmTEioCZW1fwwstaQv67RsV+t4JFh9jJ5eNf598PU6zdkxLZXQ9GMkkMQCVV0GtoBH3p3KiM32K
bWnEwexXCviRtl3wmhkMTdPolssw2kcnPLTLkmU/fY9Um+trcaxPdpDck14+5jwbbMOqgCBPz/dN
SwlnzlFG+oHdMv7bIQ9RJcOZvYLp0fLy4TTvEZupkaXWE/xeMbthK0fpsQxYt4bbx/m4vS6b+SZA
u2G+z3uf+FmRTMOI4jsllyrxd48EN0+fTuuu47kVW9vptf6ZkBDqaMmFBzHtBHBHJ0dCkdoTr7C1
7eKj48NxgssUa2zDt9I+BbMfyxemmZ9r1ZLENoIk252c7xwKrj3yeIwB3Lr5D18VMojALFO8V7Do
id6AjQYMJA88UwtzsVmGPQ2dT4CjqA1ZoymBd8OD+yQJB6rAbR8E/dXsZewUQCOZFVCrwbk1+QZv
AbdPyf9lMDDCkyKdMZ9XMl3+N5UCJ4ix8o94HwMh6QqUPQ9UC7YxgPS84OTyI9onUpiZUc5BpxXP
DwyFhHbpoIX4x9Y7s5B2HU5ctXp6Sk5MLzXhgl5lrEXw6hnJ2daWHYX+oaSMsIOXNNAfAdvURa5A
NDU3dce3MxS/VH/mKWJBIHljcIIsu8Fk9X/F78Jo8jfmIxuNM5XizYhjiVVjmkPuiYauYNmHoeND
lICVl4lQys3YECHELsn9Q9sNRoKoqrv/nFUd0AsUEBuxEQ4SeoHcwE2/v3foCTK+DAqIzHwaETHq
NbbolrpokX9z0uP/DxnylnVAoqt8sGSW+z+2nbqV+vidp6aY3CannL58r1E7wLvbl5pF5XZsTjKf
ILB2jM/nqb3Ya2I98Z18pSYnLKry11zH7F5WGe+mq0wvT4mLwHAFnQBZ6yqp+fWh6aXLeV8B4LJo
LLZxYRIZvAp3KG4C0Ax77lfMzZ8R3LweBoSKMnSFrZkOcx2YinWTVoBUCY90atm+E7Ap19ZhjTaN
skdqXjlZeH/zb0DIiSzNDOrGC7OF61ttzn7s8HE0GdMkS+qGatrpaksviA4zjbdY/uw1EAi+q66Q
u6/T1SqCAJZiIpUibmxPMydsHfXAf0aRH1bj4Zedn1ljUE46FfV1FWc2jBaK/jedoDEbsYdIA6Ua
CZV15an6EPraHPGRXak1/ns6ElLLpsP21TJoWpdUXhYgdZdDVGb1QflJw96WNbCGg202veNx4Om4
qQAGosiMG5UpfZIQC3rq7Rw5tJiZIJOuFa1spy982cGzDcP6+nqlbe4AWYLseBnR0ZMdE9e18Wyo
etwSXLk/8NnjwxXGKMLXUv9DdQ0PL39SIYZtVZHeiBzN2lBD0PZ7atwdJvEWYbVTs7ppqq9g3NIw
xV+r7+8mN4zjJADIj52HpTxBRGzUi9ml2DZ9APIBcbTv4VTRLjL+OhL8Cu/PtPmnXbusUOoExQiC
g1PZ/oIHLVnKZLmicOm/yhhdK1dwhQ8dk40aix/uXfIAUxjbwtzmdg7HU47fYfPgrcrAAgehHAMs
RN7ancrY+z1pRun8PeLuc9anxfktkB5Ohb9YvQpAwhXE8SdlmrZifRvT4cF/EhQvcQq8ECqFoUnn
4JWpXo9X2XNEROXDSqOUmYirCuwDyFYEE+39gC42COMkLPqn+Zh9N7nOdplcuDENcHMefWaxnlz6
9S8YEHaDdx7aYq/19+cv9D5NQLKUm+teMXOVTSlJx1a/3EIZ6ioxS2UiXAQL2gkda7GfU3D8v7lc
2tc0JuNK4QmztvvHo7cp4l4umhKk4+tjmdwjkif9XxmqlGsHN3LyOkPdg9e0C1MNR8gCkMOeOwcI
WbWUPEa1c1LAeYH1XBLu9wjWJVaG5/k9TmqL+boKfF094aQoM9Ec6cx4LUjs1E4mtXVz59kiOlE7
YkbrV3+axtTnu1c06XqrYotPUExWr8ZsUiFhpn3jTiYdzEXv9Jce3TgsoBxEFZwZQSQLrl1n+xgf
bmP247eYV9L0IC7b+B2V9MgkIkyAFfelTY4pYda8sRyg77PbB9IWHMs/BvUTWLecWSJ92ejAjGvQ
6Tlx8tXGnUdbEQLyCEEdSwgA0krwM1JWUfgm/pXX9Amowev3zp2deQOKqEpKZ0kmVJR+PIByCzKQ
Yxva9in33ZGsJIVDZTLaBRv02KIaYWP+QLt65blC3W/vqnXHvMDIAm2Y+OJ9M2I7/v8I5IGtfuzz
caiFRcPzxtVgzNI1GFXbqpy5GbGc2m5lXO8SKJgtfooZavVU6hqH4Srp6ptnbTsOEPhQKLUU4p7O
I8IssN/+Kq7A5cMPpbMkCSgzHIoedXrPGKqd0uqoxYCr5FIBbyntfQPoDCYm++FwXfC3/WuOvS/f
xD2/FABTTOgpqEeQGuXgaSHTEUw3Vzw4vB/zzQFR8yorcALOD26uC1QQWn3/W7P3+jlUF+UwbTYa
2tkAFRwtllFaW3+tA+5rjlZdA1/7VTPCo/6B/Sgv5jMxp0RtJtN7eGG7vDUtrn4PdVJ7YbuHsJMy
K7TYScXjYXq5qV+lzDfJylM09/bRFAmOVyHJSq9VyuPoiIb/VCjps76qx3MJtRWaLJmo3oRTnjOF
TlqZwt5P6Xfg/pWqjuhTPAFR9uxZROfmOxjuNymCoDJkyfHXzO9QEMiRa0cZDZyIuoZ/i5SFXxz8
2T8mSgp/69cTvzXAKfG1OScH7U77ZolYHprHqMNY6hi5haVV4e/TLB/PbpAXyBJoDW+GKjuu60LU
//8NMyQtcZs2bXrWWYadRypVBqEFelHzNE81ImLSGtC60aIvuc4BJ1sqOBcTa/6ixKx6EHyuIgpv
NN1I+kROc8pJn2T4roq8NDSWbslwwKr3KmbJHPG9+DChjauFdBeyxHEFxZz5bE+kI9tUmoJnt0lE
bXnSnt81xje8udsGd7ZJxqj0Akrh8vSqXHx4aN18tX1s3thZrHnJOzYRGcaLOA1hJUIWzZHENCHT
zvpWqRapzeLFo7SIB6QLbcG4BT/4WaeJjOD/J68+jcpVw64vQ0dcbYzPdjO0zhFHnQsOK9KSuYNi
ee/JZOBCg+xF4aNqM28UIaz9W33c7CRMpk2qWA+u+USGZtpp71Q+tl0MoJug31vkaYWdmdQUhtpr
o4wptXCDx/oOjTF/EigrKew5hwFYOXpeTfGrVMXjnmLjAyitdTjSK2HF2Q+XIlADosKga4/C03z6
dRNgAdDFn1V4iU7n4pppcWA+tvhCLLFMezPfi421s6yhI0s7vwCIpNPLWIjclytxFavKa6189DtN
BwvtpIuiSXZy4w/lYVY7pqiSPMobSyWFHplsmksL2/Xwv+JhQAvbVEx+G2FObDWjj7Wy46B00y/5
nlNhwXjz+Bir/97k7/ievdJ2NUlw0p/QQvxJAKyJrruSBXC5ecaV+sdRbVLu6WlZJ5Rx2jkN3z0f
sJWmvY31+CVK5nZSPlG0n0QjdL0BDu+v/8hapoUtfke8NCmOIDqQnJ/mlg7oJ/mRBTa7LyDkZIkq
T2/cTWh9YMcL1aA8kt/V2Np/8rAKTzvd7lCChxnHodvose/4CwJwUMmE24bJsfiFEXPYWcOKeKHp
wGcupITcu8CzzXOkKWnaOFVytQakqEs3k6OzZNJwb/Noj9/AXM8UoP31AXoJzFEaJAn271rIqmtD
zkH0NzBBP2MMN1Kf5okvEnRIfhhyNv3waF3U2nyaPWeh7VPcu1E12spPFvTtvKe7a0RZUonV2gBn
h7r6O8mp8E5NdeS8337EhIRcQfNeoB6WlGECBtMlqHaH0Hd/wtj4kEpDu8wgr8mnUo43bqgtKrdJ
7n4Ku0ZcLC0mI8tCikZd27kCOBttAkFKf9wx+47iUuUPH+/0a1dGwEDkjPY1H2B9seouCLAV9fll
9a6nF+grFiCtpLf0gPYkP+1YGthxsnQQ9J/+PlaO0mWFrUJQXwHlxYRcBnSFEqe9TqWWo4H4M3H5
mOSHkhg6wfhLFMR0P9hpVAP/vmYT7WwmqOwfTmmj6RGjQjhMyO21VDaBcUZM5KGPv9KPh4hVD56m
cYXqbEyQqkL+wpPFAJ1j3R3QYvYLb+5HtFy2yKm9w0fRT6JipfXDbmjC05V4G0k369WMpSNTwL1F
C2LKEmIvCGG7lFJsDNtEDUWUvzjOoNuQVxXs5OWp83oZrRabpHtjWzb0xkXHZXvoIzTUWlEFzBem
2UI1bKu/Jvwq5yOopjAx9vL+xNUnR2gnwLV4e47yCQno6mcbPc3AF1horuWaFyVfwZBO9vumCrDY
r60Z+tvu6D6yX7HpvrVbIgNDjcclsj4kZRtlhW+dyQ0Tx9bljnawWFzLsIgmcUiPxjLKujFcsz3f
e6t8+LsdTL91aW521pAJ9fOMXIy82sTMF6ealBMrlvnxi+JsXV74HPALNhBG6F4ecYXy7qwZOVFP
6AWhlNft5eKs2BrxRIfEJ29tLs+uVB/EQM+pIH0N3UfbjtFlIkTq+SL9ATSI/OVCrhdRKQtg5cpq
LDxExWnPD7ni7/sqS/VJq3d1x0RUOoePrhE1rRPBhS5xnlGryFLoKpiSOTmTZb5LUxaTztlGVwLR
de7PALIQTeOM5ZzfzmHmg2TobKbz96mluNnFm2LkEvjEDkdLWWgHhNabYccpoXJ9UoQ2HUG5x71+
q9qaQKvMKwv/FkXyiK/gYGruwEfuKPLzEfgHa0yeB+GUbpKQRewCUrzAohaZ4JWJcUIgz3416c//
EuEEaOOfbn3OtuzLFp1pdNNGg6hlCtjxIZcpsnf6u0DOhd+Bhb+QAtGkQsl/yiOHQzdkAIXzjrtd
SuFua0d/I2vx2yHzcMY4sHO8nDSn+K+u6qSOaj06fx/eOdLd4AvWbps3hebcYRSH9SdPSbLskDld
SV7Zm9yr2YwdVvpg9dKaooDumg9S21GGw2+zqLi57MaBEKEYCe1TvATc63jn5JBsH85zhCHFT4eZ
ixHqBGPp6gi2JwFGJzfvNOtC5dtQzLcrlCDtwPm0zbvnYzliVgAY2lQEIDJjdI/LsUkkK2VTtlu7
BzV1vF4c73+hDnSNDPX6BgWsPnCDytzUg589Gxe94orIOde7GdlOXGxQ8aOWUd1nGn2leyzTwc5H
912Xvp/ziLP/H36l4rfvnWQJUIXAxs74y0tjp+IciIRJPCz3x3eM28HSIpc4IIm5TvpKc+lv61Yx
uHVoiSLBbo4e7PLh7DYF8a0QNz6bxPQosbK/meKdxKjKlLl1d0crwx2DFp0wZxijYI1cZWJoYdzn
5LHpZJCInDQaRX7haUx5DBPxrhALI8QYiuRkjYmnM+Qzu0wTAZuXrmn5VHRUxQdB4YVDNMoiXapj
QE6VilJuN8ZviE2vbdxfO+28zFRdBg/KjV7FfVxlcjILsnd6Ek+8YRroo6HNeik0fuQRoyGBJnIl
wT4obrpmz13eqcmG9GLBmBB04MsUHIkRPVrXFCliT8o5r12qghf1OsI/HkaKuiOA1Dbk1D4letrw
LclMWuzjHT3AbW0fDn4ULdEQzg9N7HQD3CdTuyxYg32L35nCpL5WJdu33MlosTKIZ/lkEg6BaOlm
TOFdfjmgRmtcuAobATxbsNNijBtxKFX2uiXIFazqnfbNAxBrGin+IuBa65AIw8ovdVp8clPoJHHK
OV0c7Wyl1pEsoMmSabl0Cvel3jjbB2OnaVNs3SCwlHEbzzs4OqoiEmIPZ7maxqP8iLF8dHnIVJLl
lubbbrfovysnM509Gp5EAD5on9KGDvlGu7qjlYVgwZp3ZPQffsjhCow4ChYZeYHhIZaJv9q/ptYU
Y8WJtT70OvLJlYJk997C8tb/ZOullALTLa8+8OYw+pJ9WhyemP5c1jRYmknDNXC1ZStWTk/3Qu57
yPcMbyujNkfRu5dFfrU2Xp7XDWq18uBP9Pe3HilysNA/zOM44KV81zZbttt4VdzwLvWZbJzYr7ff
R/j1VcgiehUafR9TWzp4BrSRD2jRb9FG/rlbsFEBqKVrquXR2W+dZ8FW5qFuuyQmjF7F4iJuLpsW
sb3SFfHZOGehs9WLGFlp7hDc4w0PMA/MZfNfEjTknvTniQ4sz0udWFcfz6ORd4ijpPNSK9L6y3EQ
UwTQp0YUaxexppPZrkLSy5jMksX8PhAARpe4Y/muvC4RUKgclzOVvvYFa58jjyKVeCI29HI2172O
G/87+WriYziF6pzvIBl2o14CHmRIyEfeKXN7RtJlh2BeNXVGICdVl/kxOzZbOV40oRKNoQzvkmgg
TaFYbYjchqgPSjRNWkca4EDCL8GtAZmva0NV6nwuo6ojKNivGqMymN4EY6FDVJ/p6+3bEQDe9LJU
w71FGnJ9Bj6xxaHXx3BxKY6IicqqhL49iXMLkb80QoGGFYv214JH24G7/rDN1O1ez9GyFg+tgNuT
EbSivtKT9jtyLJ0v3jK8oS1ZeaA2LFB18aKPCug+aMX3alrL4TZIVGE8ksU028CEsFbLD4vsqOZe
Pnyo86i8H2F6MFkJw2EVG/6llFTaXNKYgc/ixrCWZ/uUGqxlyfZMD7kMCXi1QUv4fKyzSjRj/ACd
vRHmPKJ3o6PnvGe8ENOwp7PFgiUYgsgh7mLAyZ3iz1Hg0tcxYtztKXu8knE+s/c7RYC6tM+FKJRR
DkT24f9hOb0BOFYE/BOphXNfxffePvfNNOgrA2JoP9M6FRsISXMk/x67NFyhsUK+B9KNoXyOOVmH
53XQwZ8rThecgnsxBwX7IhZ6sVf5R2F6deFRLZZ7LuJDSYieGAsu7a7DIW9DQr8jr06DBlgu2Pl6
ZuQ50gPeiKWL+sbEOdm4BGG3NEdIYBWz7V9rDvNjdqfLlvqSt2pkGPcQdekNOEujN4ZGAWZsn0uv
lg/xQrMxfDKuH6nkJ5EPKzQQUeYLSpwTMFNbMjuOLCp2U7tG1G2w/b81mX2Il2SnA0lK/LFXshuF
+hZK16hb9+OuDCVNVEMqi+UGShEtTRW2a1u8G9v+s2GlX/wEBg2kaSYWp30fFcgee5i0SNo9n8By
cET/cAvgcX9sq/tKxvqC+RLHooWMfrX7qe8FTF+qCVgFjxWgjav0tNHz+HCtUW2jf4k50kWC00O2
NQyE3QJ09F319S96j+f7TnicdVM4hjxGIRTpI/airx8f9qefiBSbTAdqEr4jsgdB87ySHxuczdXx
N/xBrM2OJNWHhXoaf1Gg6EpyHgwAHfTrvW1TGpOFA3JWdzFebet0uu5BVQxEa5CgxjBeSvTna7Bs
jL8onPLk7uABF6RKqzkgGBzRmh7tC7IgbwJawp0l59t+ndqcBOE/uA+0GezXbWbkeX2vGfCo9FbH
gbKFaqmB1UKZnUQ4RqCO2Lh8LtpVBTTx80Kjm3SGYN0HCYM0NsTvr8rkgJMwei2CX1OTE8VJfDkt
zERV/TJ6ShFQmpXHLpDSwrSoRzMNdfW1h6uNpEIb+2we5zTgJxu++F2A7eJWJIaRF/qNbkcIa9jw
Sb6isrdM+HyQeYVVFCjt69ZQfJmCMdKMeYJLFjB8m5G8kAcSnelhs3LIkODtKIQ2epugsx6tmIIy
4hDF2mZSgvy3mEvxbEsZe8dKqn+KuXNsOGEepAjmm6v3BaCcAAKh7fnCO2XPlfQLaRipZnhBfIo8
VZ2xZuBwVbVTfvIzK9qEG9Y2N/S84aYV6UmhVNyWu+JRlJC5g76Jna+XNxkmCKXfysA5hHoq2WwP
9eZgx8ECsDn5YDdhgwuvr8DtTrecgEkJwASSOxcdrrexFnNwik6SQ8TRqccKg7j/Bg55EaRzmGeQ
EntetnrHDNV3Cr5oFqZ72HC6pdotuoNDSk0DEf/To+OD4E57mdE5qeJj6gFP/JDuBXJx7FhlAu1q
9xrokCU7ggEiKHneyfgiI/gAmMNDZVxMTPXJtDGGaQhalDbn7yqX9cKidhmSL/2rinj9Pg2QlP8/
E1alqQ5KBAkwv2t/Sarhw8yJ0XOYkcxb5nHXiQCqZ7yzs5Y307rL0auxYiIZhU/l5KUpiHcD7TSK
qbfHb9n65f/kLHHilIGK8n3C2b5T4SMwcJl/7ZkmKjVF9SQa1H+D2mu5tle1djy9tZHWo69KnhuB
/DpEi5pNYkw8WFvIaxStqBkVqN8Jn0tcq5zPuVth1/sTiUtjkbRsagYSIiWWZ+OSWP56rCQ5vKBm
LbCDeZRjli9IcTnVCyKIFJumaa8snClLFXVt6UVtcfuunuoA8fykSI40A5w4ORuC7P5PgZe0xSph
PAW0AupMf44OlMhXzcxBISj40VFjrhWTwvcXq1whn8UFhrQwXptwUcesX7u8uDJJq42avr/ZK8D6
FAPtFOAdjah0Pp/sg96pFcjskVOD/NMsldW1VZmK3sIpz5BETbo1LiqdOzhFs16TY8h8bMaZoytJ
O/0VCSIU8tWN4SP7ao8t+tVVu9xyxtFpmqWKLSjWz/9X8gEm2xQZzq8d7EhGzraFMdEchJHRLv2f
XMlbeaSdWITzWM/KNmtNzwuTzcixkXFicuT0AGuXZGcTnKNJwYQFoRRCBkOTk74bjeGIwMCb0rqV
CcgZYXpI7yu0pEm2Gb9+Wy+FrNsWJJzAuTWBw/PIGxqGVdqPm1f0RAkJnZANUed2m7L1YEjDL0LD
Dvn6UJ2qt8nfkm3JwDqJ4yKILDBxdCI7FGxOxAVwWvqxWpqHDcs2mZAP+mgqplE1rmdCBHokVns3
7DSiUyZNvSrkiKY6MEuN7Q19qb9+/IA6ZcD70D0YSKxCK9z2d0LnQBZtXymxhO77/ERrPspmBwqr
hFYSulszptA4LFfmS8LtL9CvO5uQ9Rii0pPXhKw7O0UPZgUXccwegFF51/Biu34d+o/QjjkjDwFC
D0X/UojIwi974gTFvboWpOj8nBEQc5EjwYBpL8prVnBJxMj7U9F6r6Us5x/sMKU/2yHimRRFJO0o
mifIygayMTUm+S0B4sS/cSz2PSm2qKpgImvG491diEOKxRKlVu9G5ioldzE3CnE4yevL8bytklvH
m7bHMLVBWdflvHdZowjHuSwzC/fHafpaNzjlcR/gwGesfBkSLjDxIBwMjl9eFbwheR33TUqgvxQq
h5l5wQmEelkNi9uJperRzx1D3RafRv+7PZXeW+gcuXIYnUzq2PK9CDlVDNhbTMZhJIdFdkQnwAy7
eAwR8t3azcEL2p3vE7Ob+jZMa1TN8LCLd33Q+GFZYkHq81zU5cD9UgbO+aw6UyPuqWIMlT5h4P+T
xqYzxLcDM0Or0T/76O/dGJX+n1YWz0jocrgA8sqVlF+0ytMtzHoxNAyKKd+AjXC82355+7f/hXS3
nCtgoxfuSqxyD2CtukMvGCsjujWt0fuSr2NU7kin0+HHMMnWH5CgPIDHp/3ClnteHuytx4VaItEW
Y5J6vuSNWcED5l7y+fJoN70+HkaA7MY40tlCpT7p+we6/mMKYzEG4+tnNuhtDmPtTqYQ3rfYkTz4
T3kpOzjmDc6oHVo0ibHJw5hbk4xoT3ujzaeIcT5mkA30lyieYU8DMoZ1U3jFpNG4ue5HI+0AKgdb
EJ6nqyCglO+wh/3TDOECopzdQOsJbV0U2fVnrZ3JJgn9NPZCclG4YH1otUBH5S7dxvJn7FSiJKPp
BFEWY1agWIvpU1H6eEn0YgVTfWb6W99qJm86uqR1b2nAlgKAwOewPliQbLLCAArmqR5EWY7+1XFw
dsUydePjQmMkbECuMBtfabwESjsTak5PfBmR1t0XvIgIyaSZrdGIymznJpIjma7qleZKmUUzhpz5
mu6Q0UwyGC/YKSRsHmybjI1YXJiISy7LpPBg3OQGpDOa8vd9yxZ9/iOj3lxVJ6NZGOKrFCtv9qxG
l/n9AgBoSVoyzpBWEh7PxJh+yFwZtnb0Puf3ze+cjGVlhw4/qurWkQ5yJIhldsQOFiYlR2oJ6nOv
yt+osaDVMgEnqOqUIqIamezgt5X18vqGAX80KBWRrSOE5HHhZ4mAf79srJaPHP9OCUg4jYopT6ZG
HfGSGRv0zbOjjbHi39KDstWQxXdci6kAEmDZXXlzo4FRrFPpF/5C4/39n1BF384ECzgwK9QvKOv1
ypTix7hz+sSPupoXNrz1f/4soTQvtMf495IkR0KQedU0xp70d2yV2TmlezRGOeYXltFcC4vVE4xl
xBQoDqMzf+Lvo0FGB1aTjgMb1Wlo8h3vbmLTadQJdBClCbkEFifuchbO7WUAmwVDnd/cHbalrlmp
G7c1Bq318gSImRXrAe4tQ9aznUlIKJvla5f3xUuYkFh7I+aPUGIYSrgO3T/oxZOPjiOc/y+9HVIT
vb5uNoaae/+WYmvRFA0BQWBCh91kmQRKB0jJS0zHLIvac+fpwEkGS2io2fYrQvEcCrCu0hv7YTAc
e/yWVIlTyUaxsJ4UTUy4vA47zj+BkT7WOu6artGa/oudqyw8FkYNEeg16eYAuGRda7x/Z8A/6+fb
3mXkpguCMXAlLPMJSwQ2g43EJM+QuFQUyYnAsUOavtJCavIo0b3VMyyTFap4HGNSC3UUMbJpFgQb
kZ0yDGrLo6j8T6OegtoPvfboYKatrV7yvP//WzfIuLPospXkzbYuZBvoIMc5I9Z8nc9vPSlwJR0d
IfDOYKRsiSzd4L9sSExv1GQ50GNgTMZ9xpD/tflFbZwcHb/ATSPcFYzxk8Tjf25ZRiqHgU44q45Y
6oILvf3hzZC4PUIm4psTGaVssT+GI9Ygthdaaf4C2pT3ylc5M6nGRe6ruwM9TFiJ/uFl+V5Je+QH
CiKZusotok/BL617wRi1YTHwfOWfgBTIyLU9zb6LVGLfuyPOip3G5HiPhOOmao8D3IQIFBWXf4je
x0nQS6WZDnrBcB/ZpY0bRe+rsT/FGmvVq/gEHSa1eRH4aA4gzt9oTUQ4kzMpe1Qh+Ullth3CbtZ8
uxmQ+wnSW+8WgWzp7YEq1/Hz0UBCHXi5aZAktqRCHN/3j7MU4X5n4n5YBW8B/aBiNWpi5bqnVyzP
d8A6ne7QXLOl1Yglhc1KF9Lhyv38kUVYktA0Li6OyVVbYWwfYZzxB3wCIjKweXoUdfnJRwBejdSK
bhu+DPEaRgAMb35Z5ALaWz3viqORcWCiCYJ2DYaigoJ8uujgGjuhug+Pc+5PyYbHGK24ED585UU1
hXCryFgWpbOzzwckRfJb6cog853Of5+iXlxeulpZxddrVmMyh7STdpuB9z76+/FIkIIbB2qwGRRb
IpsD3E6nlLZMnDjmP20FQOBP3VhEtgZ3ghW4pBIOa+v43htBNNF4Eyay1V2BkHbUv8l8mii0TxYT
9yHgn/33ks9+fxn8IB1Ta0/V1XVBEJFC/ieQ3LdBrl6ac9uF75xN3UGiL2EdJJG2VPx0lPLALqc+
6OQ4qhP0rdXq8jpVGTtsdK9zm/ZeXlcm7ubPCS5/C2VacqLmPwyhbDMSsu3Mu4N9zMuRcqSXU+ti
JwHF3zVKbS5I/ThA4gFJKHq5xvQBzOzzvlSRSRtHX5k1wI5v208vzU+lGGlzC61p2a6v48vR/oxS
3UF6O+nrxRsWwi+tYjSwURJSoooYh9tDhKmm2H8WxqFbbnv2xegxtHQoV0o6aGHdYOpws1ISCQZv
VCy3HsZ6+DMDy1SAJ4ZO1UQ5Xi9NO42BfjrMWa6ja8rKnvCAoBICsUAJr4TQ3CvvLPEy0J4gb1Cc
sbZg+IMQyYPdZdbkz4UDManVcqL3Ji46bPC/IltnXv2ex3KeZlfeB3i+HyeCHhJ67Dc8v/FPKF3f
BsnrocxBCKCsElQvaKfL+DAp/t0dRCYLs2XWK8W6MuGFErvq4060NRjls7YQ76c71mudbgi3NI8v
0gsRSkh4bRP9w7uQdm/TJgEwZZVDl5bOcHD8uGoanq1ignzKkbJrmiT0tMHaxfuWDYsrv4e64Zm3
NgczPSDf43rtr3lIk2GWf9IefWU17BjwtanQwUKxnm1260CrBc7kZ4eY2sMVfGEdA6dGnfT67ReR
4h6SAXimf+BU13K41EEZvagGpLzRTCiLIarYVsYpSfivKrTLroGcKRMJ47zerqhA9qIN6BXqNL/7
sg0cd3gmtXHqXLUW67IeYc4SPBdr7WqaHWNf8vEBBzQ4bayb+Qg3a9nBU+EwoZr7BooNUh29rVb5
Ad1VKykb8hj0AmdUJcT2XGauaIOpU4RTv62z0Zb/lK/Kgr3/q41mWK8Cyo3pmINqs8if+O6cmb4A
opPBFZGkiTVrKK+EL33SPpWCpZuXHFNzU9yeyWPxD2e4nD+xJkV1WgofRsBDk/DJfq52B3Cvuc24
13jaxXCPLWcJYbnd0t4ShUEEtoTPMnKiVg30xvx3PdKC5ExjIswboDaPBkeEaMXxADhG3H3kd1Pj
ZpuubVL66sxRhp9RjHQsoi2oRCZ7p8lV+clcya8HshuRW6K0nD/VdLeLyMq7iV7WPW0HddfiKnSD
ufqeL/NnnD+VTFVIGREQJR9O0k6V0aAViRK9blJVHPunVuTNLHE866qyHWPJG0cvJoLlMhym8MQm
gJFCe+9FJofjW8yhiGA7dyz91Gn1IHmX6rWDeqIJ0G+7Jk2rrglysco5DG+hNxFMiVv5npbMG3sV
Jo3Ve0p11UaZ9+cTqZZK7m7v+56EcpbrBTBssQ+7/g4/YVVmcI43rnN6fwMvbxwX0JVaJkNZm+0L
97Wtwmb5MW+NcSqmbWMgc0O5sI4vWt6OvzI/rYq+p+CtP2KoJl1qpPSwiuZkl9RObR2YROe0oDTW
j4VCnl/HQB2SIMMIQL9rnxSiM4fko//4i7H/OtYuh6yUHW+egB9g+sLtzT459/YS6OFX8YAzBF9C
tTlvCMs3SRSWMrK2GrloyZgEaG/x1oM210g8YQgdN3cEqFqcgKGH7/Kfwk2g/9giVxfCoLHFrusg
9QyOd8x+eSJKfTnQOfDJanCHsHf4z9glVKDJfKU3nsUDAxD3u0KSbLZF6LGdLiNKWoFmqEpJXqQd
gY9vb+D9a69Eu0f03YZ0WRGZvGgq8M5SeOnhCXp0PGKMOJtXO/8mjllbyaUYgqPcfN8vd8qpURK7
4hU/6aim7GezXJ67+wRB3s4dmi6xZqHNjWHsEdkI7CIfZZ7xlFxUUmtWbD5/GIdLcjQb3dAh1pWa
BUgI5W/yr6zastzSbkust4cSxbMnwN4JI+9tPGPOJb5kkGowex/dxMPU4qaOmLbOGeG17f47iNt/
dmOuxXnge5hM/eit3DSdKv+/QIaMFBPHjjrABQHG6YIt+OeZGiXK/6fTCORrNF+PQuAb8v3wBG0I
/MdJ9UiHb/sYGqRpIEVRkkj0GjbnRtUQA0sLXcK8BK4ilOsnbXLjw5KvhZu7srY5D+SfqABu/rvo
jGIDdlpAD6gK1W2mE0/5Nsi7qB+SLbKh1T5s48QA9GJgMCrJYvsjWFjHtQegzcdEIas0FaGUhjQg
/AtxcRL93UdRgbY+Pu59iX5fPAW/wGLSRDFmSWw4b7PYuXutn9twp/SlWR1IZ9tMUQbdItCq9kbA
bneCivBJl05csw0+/ziiBiWRL3hBX7WVwGG3PcXuXwMZcvPXudFWstxbPyGveoxb+xvopzfuXAKI
ITqETULt8Yys1Dz7d3nUk61h/RLUq/Yg/BgiIDtmYt1pLBQlbmdJiXr9kfy/K7MFWdcqYqlhJ6/Y
KGnmDcGSjoeP229tMGr1p/8UJkUbZP72tGXNVbxoXpdmvvlc1C4L/tlqZ8/GzmNyNfCpOvIpoz43
Ng8RDJi8f2QE3+rRSA15goc5+rXnJCOcl++MlvvDwMxgHc8RJCQhGFtU+DYguMAO6hIC5L1jRBDT
v6sbWB8T8RUeX62l1J+0Oi6EE+PT/jPgSjtbh72N033QZcJAyqtrxgUbw1Xv7NBquWI5WwQRBE3D
bom9qvcwMw7nY8Sh1s5tA8emRmnyhNo6YMdJyWSkD1LaO956gi6Wz/tbYZguv8pT5HS4G2TdNQ5p
S/+EFs/xbWBDg8R/R0Ff9qtEdQYfFDCvRcmhVfGIKvcbbT7VGl0undJ/JK4wdi9Uzy7ztflrXaAo
kpAmYr/iPRb5Io95z2dAPudsLrq3LeT/sbhnNtezyADHkb75MQPyTpCTo+k73EKlJCIPDK2Fm4kX
aYGMLVktUWTQ87efnjFQTEVQbS/svAFUTtjUhWit1YVkeU1YOKuI0w8pWyyEynQlLREPiy2Xf4z/
jrvdrmHK6QlA8qcrmEX4F3x/ue/XquBOmnGx69h7v0YRWIR8a5jHLECxFSZfc4g5kX9wmKE3FADe
JSFPx5ee9nIkBhMUF4FkMNJR92OljGCzsHwNBrVDyGuFY0CY98aLD2OLXa0vJizVmlHcaKGNgegj
gB+VgKG+OH0ck4QF/Reucg76VmMja0gb8r8iismrWrGdxzdZ2MYM7alQXl/gOzMBvJqfrcbtsWhd
I99rocwDeO6PJi4Zs40poJ6kr6DIVamkAewoTtM3Nh0pPPjz6xjdPKHFVcGYeI8lvJcbcesZQxBt
QdK5YW3lxbL6D7WijMRSIku6UEDfteHokeln0lqHdsl3hSlp7ZWoiHbuKK0jMrgREz3g0L04penm
Z6LorCQGpE3S7FOMBOutS4PaXyENnu3kBml+IwQbSbK+NFDMyFyzgTVp7yN4zJ1cHbAZGSXJEnKl
enGbanQdK7Mx4eliBgLh6qsy5Q9NVx4K8Dk5YyfeUiWSMiYEJCbF8hH/+1egyfyNzTNWcqNQ4qMK
0EntzLbJZ6npx5XGykHAlnURZythDCtMYl0uzAjf8nBlzmko23G9qyAGIG7GRQWtqpM7KanEK4cD
Y3dFoT6I7jSayzsFmsvZc/TsOCUVzgFNNx7EzXCFPanKxg81r7JWLkEJfHLzIsxETBexg5ouASW0
2os9NgcnjM84L9Mci9KUPzeXEZxNj/wr/5m4THnmyAeZViPKDfR2Zh3hdOQKS9zkM9CD4Wu2x3oT
8B+nm3q7TyaSBjB1Ntg9Kk8u35xBF7ANKiwhEcrUn4eEob8TYnzCWcIsEb9CD1bXaRLSQgYao2mr
5vFE5+44TyihfWibjPgK491Ua8ydXlVdQrNo3WBOnOdMlWmRTnrK3euVanP+gyq+wjFvJwl0s1Q8
jSRhPsSuk6JEZSyazjfHkx1p5J9CN48/bEibzA+ARylw0sN4GeTEKAEBcSLqRPAuwVXOpwAgCoPY
YsdNpS25Z8FRk6+aPhH+ELV/RuEGDt7X2uFashsyBhB1GVm/IM0tLryKOZGP567dFMTFoimhmHnR
okgDvLTAk0uIoP1zgjA39mdaoROxZ90BLsKcWtkOKmPStQ7zoyB8WuUtE4oXr1oXi9kT9NG6Zo+j
49WD1vJDEGdDZXy/M73sI0hhECSSxTDkE4xHsPN0aICObjBAIY5oTZZNlT7UGL68PgDHyhSu7MNS
u4tLdHTMVlr+HelY0P4CsjuSpmZcZHCWtXhPp0vqM+Wq3++WX0pTNQeOC/KODXC+evbbo4SNi6/C
ZECaPkJgKA4hDEZnfWYaBhRjSeE1BTmzWRmucRcjaf9oOKFPNOGf0FTLO6GaG2IfxUp8Xjp/r5cb
a+tNOm/RptFyKiqKp+jc75iHi0T/TXbw5a425FPMn6FtkTQk/9p5p9jR0VAlIXpz7zwlpEBnCsl8
2BjCPOoVCGtwHCSUUokFtvwvWH7INYdgMxg51D3h5Lrr0bbKBtbwgWHwfqODyFRRR1Y208bWkiId
ZWUPo/eSvoTmRSKnOI3FR/20boY9qsJYgtXJLVuhb5s37lbb2na6mVZIkwuNB8GPh+V1mGUWZjfR
ORi3SHpt6wlr4JkZ2PD/B4PeLNjzcQdfxfiCbQnc/pIgUC+YpG7G1tvHQ+ON3zC2GVFj/hzFR5ue
tAO5dR7Y7N/U4GliX8IoLMg4biCF1gBb8Znee3xVeYvQof5MYBYI0oWF8vgR6geyj0YEb1p5Qlvo
NpeucGkGPMc8vITcgg9uEl1WxSyIf0vwHnMSAy6J/VAAsGTQ662Dm2H1E3AzNMJMjjTsIEZ6R5Cy
qJXR8joHTUaS/GtEqgNHe/BCNAgY4YBbK/3N0AQlQJxNAhUUlFVhGFC2Z/wH0KkO92BwQgvvB59+
XZ85Qqa0wBnKMDqx/BlD/ckdeYQ+kUqMVlw7lIBMD7hWZ1x9g4eQPuU+rwHnE/18u+RrfMlFiOjl
kl2CQ48RnzuF52cPwSbhEOGPlripndVr5TF7H3CyLSyZFV2FdoQc5GRjQKe5WlK9ILfltFSm4NzC
/hH3khcw9Y9UgHhyczsKxZoMlIFZSKaA4U2KZ/RMRzkyoMhOT/tjmdlWQOWgRK496rV/JIBuYoM/
oQ9TNYYGZgjlva6e88SKF6XqpDlf0DBD4usGzORLOhNdq7YcCsIqjDHGJJTHi7S9XMxcnPtFH9vO
d8uCV9DpJ+mRHhF9DbXg1sLP1XOh1i7d7nuzwLKML7QVg0Ni1hStSytPKFmZMxqLQpFoH/AjCp11
d8wcXj5GfD0FGsOiJq44Eaa5QCtllGcwyJ0AOz3cOUK+T5gxVvQ9kys0+QsolaaW7Dv6+0hKWDGI
Dl6qs+o+DjnsQ+Ea+MdIOliBd/vz3pBnd/QmncHg1HhLPgD6AJ/V3AB/pGp5ZsANpVMxBCo1ytqX
hFP7mcXRy2pn9meePnhIJa4Lo5weKxcHjQgwlkeKHZM/TA+30YoRqfqBzYD22kS16crBcCbrJm+q
ESJIQs/cX/w5ARPUaCHIjEV5BX30jKNrpD5GFrPrSouXH8oHPafBdEDbW6fA2uBQdPS3neZIvYs9
ojVbEdiGXTTagaZ741AUH0mAoXGyIjdQACM+UM6grGcmPUDZwCkFMdS+1kgJl8BTgU+5yxO3RYqz
SHhR9mFt6Ofdec3A79y6OdtAYid1Cy5/kB+edm3pBKMcdFskXgU8iMVTvg+b+VxylOVEtcgIFe/L
jvoK25kUmOOmeiNUyyHq+I8qSG/mh7lkcUX4J/AeOm1HX5u/dCyLlJxm5DSWWZR7Ao75ypjEOvgJ
HP0G0l8bNWyMaDI/kiXpY3ILEfHyRTkXl1wJOnMlWCWuGHhd85tAe6Wb4lM+iuSl5kHfJqlRisdh
u/O/9APKfis6AFtfqmZcZaLKhfci041XeShiaQmkjUtyP0WJal6qCwXuACT1T9J2gROyh7eQrQnZ
n3yt6j1ZW/W34sxOCKQJZwslfblV39QooKgFualUoPdg7JmJruMpjGbkICumcpPMvs/HKestq4Y3
hwO6h55oLFQ3/MaDHpGqPill1yMpoIjCFx/ia9+A+sGEwOXkTTK01wCKnLr774hj83/HSZsUnCLZ
w4n36VZQiMhOZ0VFxazI9RJa1MGaM9QnTEbchOaK1DP+L24sreBqrITQdGwHDtsByGYDIfEv6vyQ
s0tvRr8zonk7oYj7Q6KI5X/FUxHJaA8wJfXupvGzq6m1ihGLwMJImOMjbkZ9GSUXFDtqKJSQ352Y
kAQlqE1c+efQYhjR6OhPyCOAB1e6aeKD+Usod+UgkaixrBsf6LQpLCvcox1Kv1019Xi2UtJxDAaa
fY+bBtsURC4CgnAhSzs+CC2ELvq2Gk6kFQ4JctsHBewV1cmaNWGGNg3S92TGze73tyStay2xiyrK
mpNhqMGjR8kUNKtG7maO/wD/cCOznhgJozYrq8yTNdqUfDbakdYAnNiwbXLLkK/e4Uxq7mkHF0WO
XJi4NBVaTiJlI1p9cVJ1v2h3hgnL/wqvxcYKprIq/CZjxgjJa7Rs5kM7wn1+33um/+kuAK6DkEcm
gZDoOR9bDuBocNbwZ9kCUxpizSruAXm95OQDuVYm45r+i/q5/I/SVnrg//FKTKDJyuslcOexpsJZ
SnnB64oygkPb5/U089KQNo+EuWtc2vJYVgHO28cgOJSvabsCYIg5r+uQLe0wmmkTfsPU6yPItIfC
2uYmapxcD2o5jC8NTUpJETVyxB8i+XDrYnU1KMe/iNbcI9slg3+Kj7otxEU49WQDKJ1V4dwPPN8n
q7CtxUxxRUHBsUiphFlDKvJNCMMPmEn1i4GD6DGnQMnYaUWmbIqXIQpB1x5e2HwBXbgid74DuC6a
HD7zdFOXLCQds7+BInFgDzT4bM99K60n/dOjCWvuJzvVGrBRTP99//cjQkGaujKqfdkUJ5h+41ix
8R5aBChOm6KWuD9UVl97jsfOisuBebsSWEct0LGXgTPGM3KaAuf6h/gLDL452+FmRAYrg2VrLxER
eYn6ZxqdeiOpUeVPRkRKJJOvWt2LBX292Ncayrjq9Esg0iafGs9EMEUVnDlqTEwU9QN2DktYERzP
lQK6aKWBUt3DlPb+7VzTFH7IaC7GivYKkcdNUOq70FjuYMECSTu/2Tc+HGYHv8NFMsSPeIx0uaq0
bERfdzmE4MYEdymG7j9S2wnlnIlBamMHbak00tvn1qbtO92e7RIJXPD1Co53cos4NZoroDccU93h
7qLP4WaMsYRB26Pic8Kaf1XWLgHpsWNapgp537W7xEi2skYdNSL80EfhIfL5Rd6vPlswovt1lpiD
AUOPUpvdG/3PnxukTKypkChPn3W7bMiiR8J/skLRwJ7db2LE94kmID94Kn7vjFqz4smMdtViOPM8
0DaT5wvFI3h3f245PJ36jic7LtbOgQ3OPPjNE6j57vmSrjYjmW+zXg9151C39+q53zTAO9RQIJZg
GOHPhAK+or5FJGv8+RZO39gB5fZyw5UP4qmA+fF6CM4klaZsYAZyejFBZgJ33uj2kZ6s3fFNYrHB
o5WtEq/XPOl83O9GUtENzOUw0E8LY8TZCxTX/P4WZ9wfZgHqQ5D+TE5b3XfkRLvJpfPhlC6tVeda
4MEKKCTHdUlMB5feU8eRxIN8P4eErXNdQeW6U4iOFbZuB+31yZozW7S8uuNJ0pdyGuqQfB584ohG
MTy6ZCvo0PvcHV+Wd44zZeunSWpIipvknpatOud4hJo7N/EhD5FuKvMFHUaU1tjBYFRFT4Z/Kt1g
nVrnKhXwEss0iCTdL4Pedh+EjNEZuyX1oHvr6CSncpoI/i1oF5e1f+D82nMOkHWTOlK8qCUyWyhR
b2wz/Z4dCI2WFeiJqR7d8s8xvhWmoD8/tp7Ls0KtBmhslV+KRl0hYv8k3hU7i0uepeXJnQxwlsYH
GYpSY0c3I/ekX1Tohg5mt084+qAHzemuxLze6Ef7R8AKhupYapOVWPsxnRdDP82+OE/1Rv532qM6
6RjqG+3rmvj6erhmDAaFiiifNS+HmAndFhE33Tv5GDLOk77AYP2n5a8UL5kmRhlyuha0woZtx8su
HQhC98ndyn3ViZzYgjJoaLVv8uu54WfM3MaXbBWHnWCGY2OBLC7c9vmjB5s5MdlCgx23KczWImm9
ZyviyEo7zT14tsLZvNBhQa9kDWCVmIcFjGLLA5GgZkegthyKKhg2yAZzGQI0WZDYBKDpV3tsqs5d
oD1jRzkkGiPeZHuniSz1eMYG4wgOBSmHOvncwg/dkv38gfnWp2FTlcooe7mLxK/kBh8c5z1erSHq
gzBzhaQVGlRxltRGmvh3A9Kn8kD9JEwzd0uOqPom51pldAfJSbVBfaHu8c90BvGaBO52oQX4en6X
zkdBpoPSkv/IJri9ME1QFg9KJNIJ1+7kTAgEMIUvsL+FaemjSCdVba7Eu+r35y41CzmVmOJQpwqo
GjZ7LGrOhnvZKKypUi6n3UZ1Gl0yZc0bq7anujX01cYN/+ajgXr30vq6hzh6FxeGE5vp+Wq8/7kA
RgvTPtBRTFj9QtzMeEURnrRPJ+4+Ha56O5JGFDK3MW6pqGpCGgYFcQvkpRcvTj/ih9QaSSZ282jz
lpqgWqj4dS6yC+0ooN9izuxKCHR+ZNWkXfzJQV5Hp8GmCIl+2T8nvtMV17aksYSASJQsKopr5BXv
PmrFeoRip49jx6NAq4V87qGT+j8LRhNrljpXAWwLDD22foxHyXUeZTchTKZjxyouQEY+uzKnHS21
uY3DKqtE3EkWjKEoqEpyd1UrR0HNkib58uLVBYgM1cby5qWjJU2cpdLq71SjQIUcqwb5wvLam1Ap
ontSr+3pHm7GBWtI2rG/awpzkKfiTBN1kd05TzJyx0TDo0fIPfHr6viOcWJI/v9d5LhghOKHk+5N
91TvwLbSG24CWBEhVMXq91o9Tak1zowiMUZAzIOGfhmtF+6zw+VymqaCpFTpRT7IjH29cQB68sQX
6Bd1VJkRxYZtVDpXAj2uO3FHtymKuWGHpjMcqwyvLdQAvHQk73QAKLZAii+/oI5USwA8fA0Qk0nz
+aMhBdJljeySAnR6wkCwx/fr37UBJGoP80gZXWurRnmblArajJRs6STkToYK4FVyPyXg4OJyD0e9
Qn1GZXhI8cCrIZfT+Xq2m7tyOO7m5OYSSgrBRb/h6te5P1Fx2kZrvk3dvyAYyFAemD8B9IG3uKGF
h+royZ5SS69PTMxgnoVH9O/SdKLOtiSNIt/0a1fFz+9jrhN4en/n9x6R8UeUP9RoCah/e7vrQz71
MfcHebh8ZNK+lKHnNcf6y72dVTkVPdr/IXUERC1tEEXa3EYNjWN2rSH4SGk3u+zS5Y4WvzP24ctV
vFswJaBF3iHvuXDmxq6H8oUF5tVMd7Xziz5laIhYmbMpTVm5xrmLlingeoj6lOqDi66/+u4Kw3mz
cmtf9/+HpTJq0Lzswm0qIifzEfPXVldqO8688VP694Qjvme93xEx5m6HLKjhlxo/xGhYFAuo2mb/
pWHVuCEuoLqk76u2HrhMTQsDjfVisoCyYh+kt+mQ4BWIgL4qtkWkc0nx1tTKaebIORi14WREhIrg
zBlbJER1FX1b43KD8QRSdqcIBTPUsiA1IJUiHOQnJ3LCjm/0QhRZmAIoEniHnL7OhioQwgpQRVOu
K90yDoVjbfBN2kj9Y5d+9FHtXRtPjjOWONSu+3uBUEd3+WysYvoJcqULMm9vsp2qqIkc7fikz6/K
zgYMQWM8xWdQo0VHQFVBqHyuoBwaYZVCK0ULXIbYtqauqnIgqkElmi0T0OTg/qJXSBlEKPODSGIK
Vl937TTsNzUXUAV8m2Qz92pSHQrGn7tWOpV++iq+HrbesWc6dnAHj6aO4di/ZexMHqhokDXVpg9U
O1UdEfJe4pZgKPXvLED4qjVIL4R5JovlAtnwqabaj5QcGjcecmDpWkHjk1N0iYqdzdE+C2JVb27U
DsTXntA3oFhaBwyXGP6ktDIr2L4qTg99nByNNsk2t6I6qsca37NJEwe6JX6LLL+lE1CsEfj3Ru3C
45zmmtcNR+z/Bpr9eb2JCuDJlxBD6Z0OLaW/wsRfQJTqUHA70FR6DVqFOFfmmXqQS0L31R6co84g
iF7ff54T0N71GAZ4tMeIXu+5XXqHpJm0o72U80+UjcXEZMyr/8OIF5QWY8mObUZUg4Mi7TQ2UDvg
2c0jbYDZWZtbQh5JOMEwY9OQO4fOdAj5fu5AIJFehzpAa4/UGTADhySnbZtvKNn3FrS7n1c4GhRJ
g6ZnEyaPE0cba8SspRo6rA2mFxSCa+pwcmlUeapVWfJiIMCws+Ttykyp7p54y1KouThbVpSua4Mb
99magzpPSVBlHMp1MM9hpOP36256p/ACAOufAKfQvjnDwl8YYaFyPHqPsAKtKmC3iWad0u6IzEZa
85YZDxAuOZbQx9u9iXS0duZJv2vpZIWjuOii5phO5c9YccuDyRqSt2rJwqYfwOFzxJRv/zr3NrwU
2QNNm2J4nJkFeh5ScRl7WmYANduvaKL2P3WbDaX8nErwhrZ2zvns3byP6rEDwn6WPDJ4u9fcDHPs
65bCK35gxsU4CIGRFaeFXj0tdjyI8fHHygQAvwJf/AmZ7tcIr/VFz9S09mFa7u3c8Nv8q3xVN8zm
jS34KYf0q33fvE7zrn6TU9UoRdrSVhW65guZOhtpWTATUdaWHtSnS/owHMZtSfT3Wql7S4C80nrh
l9WTSsg5XMY0XN1X7FnErqbxKDCLVvk+OH0Yvc3MacbuUj1QlKTQ6cvfMh5YHHYAcRm4GdenCmIW
bES5Bc1UmZd0ejQMTSSMURTj/IbegsNf/R9fk28GUW8KJtyfYpGZ/bJoZjk77sNGEnHuaSeMot+S
pfBQ7BXoO/+vUFudL+W6/29IYEm73/D1whO9MPjGH0VG9OQhy6WeTuXJ/MtJctRdPt6ULRdfDoTP
nyDn0D5/BsyGAnE8X3cj2h6ewM93yEopd5MbiiFJT+TFW43E2EtoLXY67mCOWQ97y4F0vGzEjBUU
0g4zfzomKTpZU31PpWeuTXlywA1Qm62w0pd27Zgse9WCueSmth9lEw+EsOdgn+tXGH98GPPSWIFU
RKNIUwoTOI5mAATooR4uPrsoozsIulKfIgR4nQZEf1dr9DO557DlMF1XDaSMdujgWBW+d26JYRp4
Z0wwhto8kFF17JV+ommSiwE+ylXJewL0HAKUkFEX4t5JCNbDen8/8B6O/KdXbjKI6IoVILCRNeG1
i8JqFAwLCz06COGIyyhbtYPZcHNW2W6pAHEovCAjnNKJtiSsQBhULu2pr1TMHBgxKF6A0T7QMHAQ
hjxz3DLO4YEwswLv27ovpMcjzsQnUtnQoW/j6AIqS+hljOduQ6JUNUPYZkoRRFBKsiti4+EcDrxL
E8C1qtyqvRWStH75lQhW7p5kkCn1xCNEPCZDK7G98Juvd356hcjCLtB9rVKqTI2Na5cj3+vfOV+w
am82w/O+b6ii7/HVcKT/k2wuKMXj06E6yh5gzANf17TWfFRbafqfJfCI6O0B6NZrBWUAXceifrJ6
N6JIZgyb2x5vKLOeAxZSu4OIXN+Ivut0Nj6b8chv6jK0QhaOAmaWlB3urd1JJdFdmRfawlhbKOKc
83+p4ewJILfuVk5H8maxz2ube2g5/ekxvZcWfM6nXWjmK1pfal895Z0IzC3zJcOGeahq4m2IJiUr
p2YNrzVfqEH2fVHEn3j6qBTfgVunhqAIXJIIJm3La6HOcl+GoREo4AGlyLCBC9RiAVkpvqYkSKVM
N3ld2us9tDXuhkoKWjGEqVDgmXk/gy4FmE0v6dnSoXdXlL15+wQj7wgOoMYoIwsii889OrE8njGW
yfIFkuAFYMoq7XK9pmAfEUjWbenoAbEaZLxnSF3xSNrVf7Kv8rL/Xp56emkNZYDaZgprAYP3vPF2
cIhW6l31jFABPfcJNgXMB/DKkqV2bQpUCdB3zmMnAE0bda1R8zMaarcwx4Z7hmCARS81g94KFfzG
ML7A2SiNN4/MO4uIsuGeqJORGcRwWwSKnydzLkNOlN4bM5BfYEWjdehA7o/lYq21IHkHPAL6eqOq
jbcuWmj86hehX5qXppZknY0Skn4oHfTv0KRejo9IoQt87AgJUl/SSXLU2wo7YaGMtlsBFjO1VP+E
qS57mh/VrbRsJitXF1z79JAO2xOhsshwHohYQOsz1gQv/YCeg+kkXNQ3JARZI9+Zp7+fNAwa99nY
iv46jZyuK9cMXVDVJZSEG85H3SNqfg2NK1oXPCYNN9+6Vcju5+8rGF6pTA/tB8A84gkQm2UpOd0j
p45qw3PHGu3uXs1SINEPtsZipnhmh0RT6xUHGA+qECEyJ/ErvSQjCnqEYNVrwwZ9y3WOBVaLeZMU
BAVqlavPpSs8wJiADJULt/XhW0/RJQNxHVibBrXLZeiljl7KpyzDFkVfGlkvqfoftuSdeR63/NTK
NOpN3H1hfYLnGHwtTkOxFdHL+FLQIr4gk6+dP/AV+cKl+D+BY32fJ9axHsXciDcpkITChbtYyYCu
H13dF9NN6ibl4vSs4g+4ucOc4d+cLWfqENj42IHqg4xzWvbIRK2VU8USFDbyoL7bMm/i170iNxMw
l4CTIZJu31zsQSCqsbVi6DYQZHpybhjNADcLDISDOli/t2EUshqMdGuDC6PK5HFA6I+DspySoCeO
lVHJiK4/uI6oD8bbX3iDVpKQtSR71r5ZMf+b8vcWhDfyy6isoGP9hgH/VhyiAokzmzDlvKD3x7AA
of3t0COmlfPPuSrBIzyXufCpV/4BKTFdqwAYzEX6W6GO/AL/W90/1kU5IZ127WAqrmOG7s77KvLI
ZemI05CSzCkMHjw0B651ZFPqHxH59ZSj82p+dtpPpp0bRAGhpSMXWTt/RzGGHMrPE6FIx5jfofHx
skwQmJ5zD+j/7g17biceW4+JUR7hVn+kbvVt18VZVly4oRuGzfhWn5lEW63nAHsYxDyZqq/85F0c
n/cATVs8XNMeu3To+B5I5kkTPz1L04ggAXi6PQVcD5IM5z6vYjh2tuAk8O4toMBmCINNGJV9oQdj
bLxJzKA5sQRy7gHq8V3Rw06CB2Yq/2D4zQBtyDlotI/GvLr4xtX4fFvggnZ+Bektn6pm0dTwaOLe
pfxpH1HM6O399oUnwTTx4PFTvvsS05DTBOD7r6KcHaMbB6FEheTt6W+abGXwwtnR+MfsZtLCglie
BZ7pOkDYxadd96mPJDXd2YVB6KQhV9hQ0gngwZst6HpvTFbEy4/13NaIQGl2mt/u5YChE+Ud1zuv
YMx6hAQWKXI8plYr6wn8F6MnMMm/zkE7cLLY+jNuckZRlYMD0jrct3/2KNwTLCyF8YGH1sw2VfN/
/Pdqd21LEb15mYdvo8C5U11v2ooje8UiL/ucZ5ajD2mbaG/0v8kyGogrIqKPhPIsQm7fIs25+i5C
CgMBuNEtrC40UE2E3zjAzbMoI9OrQIOcS9JhIWBx9hdEFDD8ipMKBnFoGN3WoKu6GCcOH876XzhN
tTc1Xog8l6W2bVXO5w/I1uY3k7pp7fJHVAQMqXLWO3YzFICC9wtjvgZjAVXTNJichq7ylIp+jTzs
2j7tzgiEVtgyz0DSX4yXhmxbxi44iDmZ/T8c0V5Lq5CkuTaJ4eQ1ifRhKeugTGFMlwA8tA+XzhJd
pBBso9eLTo4RRz4Z62MWq1Ptopx9UGzAEAwTqIXH0irD9XA43IQneFv5d/IP0XTT1/6kzmzMua0w
4p6n0sI2JxKaCjaydEo9hMKKKn36neHUWeLHrY/wg7G1Iv2WeDjXhOTrQinzP0CB/sDdazii9LD5
xZb7GhQ34kBqlUID6iKGTFdT2Izq+KNzeIx9/wiQROc7QlDh9X1a+rCCZmeTGims0/3p4G3Ghp0V
4ZxgYeOCeuCe5J0yJtqWUrcFiVycV4nYJe9sYDigesrwKsCR7O3wcoRrvivPsEjppd5CStl0OK7e
0Mofh5u5Q3Oayx4sXjWxHK4ml8l2GpOedky1URNgz+d7W495u6XasdaPtKe1D2FuDgjYKHik4DHJ
5Ewe6eDAvdgToAdHJIRk07tEtRiR06Wt90yfFQd6DM6ind1vCGUe5tDPuG24Qe76nzJsUn+j/fLk
5nOTUzfPFNiNxEgy7H7wd34LQL/d3oR2WQDHxeAPvBxMNAcVhIuqSAamheB7XfFWhMDCh1sucXPm
TzzcpWGT1N9POVyjZLRCJRoLNH3AhN2ZVxRpevcQjJXquSp/jupQPmNFX45DXtEIBleZnxUThaww
bOZ1v+rBUbRqaLOsDQJsyxK/f2BQRKxtEHG2GPOD92M2db1eHAORzHlLSAfNW7xXEEoT3YTZXqi1
UYCpGCPz7YlE+AzbROh3M5chdM3cHImc3iSF524hKooKNTz5Ot656psKH/9dNoE6sAPhyGcbzOn0
ur7CuKpNHpAaK5vRbnCQIUM/h2tp+atJgJ+37gh4PDwMeg+ZdhUv0+Ve5KL9Z0FEoElS05j9vsNA
7l5oAk/PVgHtvjnI68ZV8j8viPPYhejxCeu7BjlzV2XtdG2tuivXUegbJqEbMzz6EUzPIijlWbxe
f6W6MmrXJDcexeCdWZVV/RFityZ8VrJG9NnBKzToIz706agbpHe9/w1AbQfKpT2Qkhs8kyxBoy5Y
QkwjCCADN5v4FV0+0d4d1AzmyJtP42gpVYypfdc6zdj4i+s/vkvpvav1oDn6QnKUynzEzMuYbIUA
up1LeKOYHV2I4TJ8F1pXzxPJObxbuzJntwiJEX3+Bu6H8Xh7c5er87bv6BwDe3Tm385JvXmVUrjq
hzdXY1AiKNWhKt6UbugD1ttB9Pm+sZcMnTF+CyFT9+AzwjAyJbtjoBeLUtd4eGrxsWNqZUMuEou/
OIJ7TCKQQNAM0TXRXZAN6ifjQQ5/Odis+qoFio2D3HdZTLpj++dovKYtoDZPTH37jfUCQvCg/7pB
4hKayrSPUWxZk4arnDMGkx1UzhPxj1unCCFG3eNhIp6oeK5wK+WPRw0D6LSJGXMHuqO08MVW0WaN
fPH6RvchVA6m5IvU6AA4k/Igr99DzaqI8iMGZDka0cKN+K572x1tA9bZRiJXjO8AKyHDU/ReYGJm
5lCsBr6Vj1nwqo69Za4y9/wCtdgLUOnCikcuGUfFUS5ycvEKfdGMmt+r1SpayEXndcsmoxZRpPyI
4wYvXKQYaiKIQ/3Uzb5fL+kmX1nMhk7L8ijaaAcT+QLXkMiNDMFCfoKuNfXJNRVb/LpD7dXNBtw0
mYtaxkaDKbbeO1znoTEZXY51OjJ8/uYJPzWYny9mvlynE8m/3RgNOXBEKsJHf7h2dYAgxaxc4gDN
9TWd0dednXnYaYZATxWaZN2jizx3ZPaiY4NeVWpphxrxc1mYJ5QMN8QJlobsGKMwDHDEHZYRaMuI
NLm3Oz/nWP5+oC+j7jMPE2CgxzPOrNl2Vei2TDix8nNIuaPz5qAZaqLe8o1QBowtj/gqWj+zx3rm
CwK3wgSFK38UpcQSuRihKYFZHua1q/4axyPGaY6lfvmNZ3zp+rQCXLsg2Oj7he2pqKz6Bx13aQ9S
s0u/c62Ccj/Bz5RQ5k8Ht3Cjk/OzmsrkCPVm/aYSgw9ZPF59ITgwPB1UDKKnZrjL0tl6GxrfWF3W
c3at0wFsILeOCRmQfWDco6+htXmvbB4cIxrov0bHpaupFCA06v7MP/hvvkzj6RJT1O0bHi8ZSQ2G
76LLGP03LlBIo7RVMGOdZrlBsPsi2SYOIQlz0X/F4EC+fPUa0fzENb+uGW/MlXGyVzDIRROEbBOQ
y5c5nURUKASlFpyEYYW6VbuyWYBPrM3YvoXsGx+/mdGC3P8rmMOGyes82iMcl8lpJjLVi/e0YZtc
jMZdLW9InG+9L2hxDnRl7WzZiBjsKY5UAu7eftwmOEr/kks6q9XEcVgIqlm5auG40E2DLE0u5Fqw
OUK9ITs6T/4hHKIKqw62DSB9SVgFDOa9ShU6LgGCjvWCxCO4SwEzxMape8XjHnAYkVYoM7nFP1+U
6TKA1YPWnfgmPR29OyknCvVrqsWNj1ptgS9e6Frsx/aghOZQj8ekdYy7ad3riQSYVD+lkwLt9k3l
iuPbzKzFCJ1R7Pgr/rw0rPJAJTVkprMfP5+7gFdQD2TeYRPW6EHVpmZisPDzADh0Ud1NrsmWT8Hu
4A4qCAArCIU5DeGINk8MT/HEfeQlFYfUY6oljS+8Kgt+pxY9Waq4O1jaLNnfvE0SJ7WsvZDITjtT
3QgnRnZl0W5pWqvzuKDWlnADg8JeXngq2Ci6V9VWT5RLUGmRd68m9jpA/80EMx/FRhxx0N7KdMq+
w6nbgRzBect3abQcFGqYzFFF0axIwxjUQLO6OfNVDa5Ilu00qDgRWqqFeBrfzZDWvgRd5BVYl6C3
oA9w/ULcRkU7rCL4QNbzidwWjBCN31Vml0pbh0NZAX4vFF4n9+cZaWEQmUrZhY1p43cMJaPZDH7Q
S6mcbBCGfGySTsFqhgmXQ9Yr76AbP+flbU3m1ZuzNRPJAgv0g/MUKB2uCWBWYH+teR7I37+yYi0M
wHIv2V59YP0oCeE6x2jSSgTKe93prAm/DV2wyNIaFy89NBYh5dJeIHEu9eQ0qJR+bUtAQZdqa4dY
IGrPBpsKyg/L/W0gPolVgSGTwY5w+bAl6oOcb3AjpFRXmYexXWHAfiy8u234gpatyXtruvN0xB1A
W61nXyVsvI8ihzqz7OWw4UAmI5zN31878A5YLyK38baxhuixsQUxzxcidWeEhIlyoqDRx3LnkMVo
BR2IZJYfvnPtje4hOly1wPCXHlDYiMWj90AFm5ieGTzSzBx2oJrKr2Zo7/urzdGFQLzwGsA56JM6
FI7x/EIpdNa+nFhKZTF+YwsgvMlzxGvQ1fwXSIOBn/lsxkU6ZURSXulV3x37dOnUuONmTk+41xst
R8wfsAf2XpnDJu0hio5LV61v4xmKY0UINAyVhyAiWZKK7LSxZh02jT8UR7NUAp84P0w+ldM1wbbu
SmjSQXAfrAdsxbTz/qvqzrtzhd+LICbZ2/zSTKwoZuF/yhc/cGMQOGvk40YxXGlSJH0S/YJg2POr
Fc6FyVdck/EWVvSGDKxfVm1OhM6h390LpB0JxrER8YAyzIRQ46ZVQ7JbCrR3c3Nrt1EJn63waHhe
iCtGhBWPZ8qwmlMFFDENyxGTHJ1LCFpuVKI6wDLql/5Ny81JB7pJttgAHd4pK5zZPKLMCOGTQWN/
sOc+S00YMyTB9uV0aBdE6WtxiWh90pvw7mO6nQGXFOZ9KbvIgVn7VbhOpS3HtcVP5hE1JDkcR9sD
iQLht/+RmxY+UYmMphO+VquFO9b+FKKLwnEls5KKvAwMgrlMYgwFhSVsDzPpuDzkpI1xlWf1s++y
0cdpOIP+BKphvz0d0+TYAxP1sx9wH5GBzwc7k9xpO5EWqJQ9WAqiw1cINwkSf1NWnRe3qLb5iRkK
lFxtCwOOqrt6YkQWO4QzBAUCSi1b3CxLlwxFDnK4PNheIKAOG50XyP94OVte2xRMXviPfm/yqmPV
QUZ4VLVT6DjHQMrl8eUi4Bh4w2ZVSLqZrZBy6ey3pifLTwkSXICbaUTzFr7GI/tyuGrk5m3+EdeW
Rc5BNPypj90chGMn2Vazj5gw9bcLsYYcL5GXEtfIrLPS5ZgITa/47kzApkHH2NP3WZZk9Ky0F5af
nINLpaTj2ZvieRoyFwB1FaD54WGBndH42uND5hW/MqEaDVITQqHIYqoSoZIBXKlm1ljxD6il8u+T
1PH4lx03r2hUIwQsDespbsNvNptdV43lL6OHzZU2oIp/cclJWNisNFXiV1GZ4a7+C5syrfK6yw6V
s/YjIcY8EQxaWvGRTyEaV/Y4ZiDpsvjLWlNy0ZRg5YnIQNRGcuEIQM2Pu2cEH/3Wir1zqLBSRnqd
iw3QXqjLKLUxqgSp+khs798Oiekx9uuonKd/mN2l0mwQwwmbbiVEpvOTX36ILCk02TjxSkMVBZXL
bjWtfqtn07fS7d1gGHQudQxWJBX4zym5o46ZeJLcZFiSkeYORQ5HMIe5WXeZjHihRzKaZMefSKTF
bFqzuWMdDmEnNXnjlDQCXBsoHS3+w2kE86rUmzBvaLPvWDHzvqQkf2WndbcBt5EzW6+IJrYslPBq
8+8fVaiCLjAYJPZKLCiVD8uptYn8lXrHXsFZbvdSlPQZ8MyLH1xP/MC7Gog1CkJVOXG1BfTS9kA5
wVlOWIhr9uY4y4dp8gBC34emgMvBLr7GvNo1ndJUNuShz94FvTzXcIDqwGT7+c10p6i0fW+3yls4
2bVmPiBaLL5ESnoBA/Radar67nCU7xuUd2jUeyYibTD9rFcR7gH29VjkY/pj+3SBKp3HwSLPZtQK
SPxJFogjuDH3vaFdnFbgYCLCgGbOtwnRUwrjOd4dpYN+dqtnmaB06Wkg1b8FrqId+Cd00jZe3rKq
Z6w9ldsRKbpPol/CdwbCGpJ8tCwSd0tUFIKsDAdTiIGSMi2BRzPLc166kHxbLM2cMqTkhxlMS2xg
KjDnLGFObJ66cOr1xAdytTOr9mZAEhY6HPvf5YiN3tPjZ/VAWN/ORkQteO9AQMXtVKgp49+BUiMu
wdtInGlk4O4stdjGiDH9dxeb7BcUQa7SOInncfebi2C+AmW4eI0D8a39WTVHnNfORFgZfz5bagaj
p/bgr5/Qi/8ZEBh0/vVx9VGmCCYJFaLA+d80AF6SLPDLAp5EYnfYp5z9O9dlSb4CufaY1/KG6T+8
EVo+ih3wE+Jwz+PG3+mQm/3aAPYChpp7uZZ2Na28zILVeWGuQwQ0EGtsc2fmmJfjNDg4959BOAcE
gEozDJR8FQLmHuyjPDFo7SwQKeL1atwlFmaLxUmAZZmmexnq9pm6fAh+fCgvhS/fRwb5LGpH3+F1
r0fNM8P/ixD1mmXP/xMILezUT3x1aUlKXjPhhy2HEmUQzdl6cyiewvmOMMPqVNBRub7gcmmmyv7X
UHMK3fv5ZNcEAqMMC/3mvlalOLZEGIB8c1nEoqIwCIgrQa73m1rcerpUAEZz3ZRGxJmcK27L4IUB
W6zl/KCY+DmLhlKcJ0HcIZJFLAiPlGL1odw4dtH44QWAL4CxHGcB4z9IVEaW08u8HXSnx2duXvxR
Ig==
`protect end_protected


